

cdl_package OROPKG_OS_LXRT {
    display "OS Abstraction Layer RTAI/LXRT"
    description "
Use this package if you want to compile 
Orocos for RTAI Realtime Userspace. It has
support for all packages used in Orocos."

    requires OROPKG_SUPPORT_RTAI

    include_dir os
    parent OROPKG_OS

    hardware

    compile MainThread.cxx
    compile fosi.c
    compile lxrtthreads.cxx

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB
    implements OROINT_OS_MAIN
    implements OROINT_OS_MAIN_THREAD
    implements OROINT_OS_LINUX_IOPERM

    define_proc {
        puts $::cdl_system_header "\#define CYGBLD_OS_TARGET_H   <pkgconf/os_lxrt.h>"
    }

    cdl_option OROSEM_OS_LXRT_CHECK {
	display "Check LXRT calls for null pointers."
	description "
Enable to check for wrongly initialised pointers
when calling an LXRT function. You can disable this
for production code."
	flavor bool
	default_value 1
    }

    cdl_option OROSEM_OS_LXRT_PERIODIC {
	display "Run RTAI Scheduler in periodic mode"
	description "
Enable to use the periodic mode of the RTAI scheduler
instead of the 'one-shot' scheduler. You need to provide
the periodic scheduler execution period in seconds (s). Leave this
disabled if unsure."
	flavor booldata
	default_value 0
	define ORODAT_OS_LXRT_PERIODIC_TICK
    }


	cdl_option ORONUM_RTAI_VERSION {
	    display "RTAI version"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor data
	    #legal_values {"2" "3"}
	    calculated { OROBLD_SUPPORT_RTAI_VERSION }
	    description "
        Select the RTAI version you are using.
Legal values are 2 and 3. This value is detected by 
the packages configure script and modifyable in
the \"Detected Support Libraries->RTAI Installation\" 
package."
	}

	cdl_option OROBLD_OS_EXTRA_CFLAGS {
	    display "RTAI Include Directory"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor data
	    no_define
	    define -format="\\\"%s\/include\/config.h\\\"" ORO_RTAI_CONFIG
	    calculated { "-I".OROBLD_SUPPORT_RTAI_DIR."/include -I".OROBLD_SUPPORT_RTAI_LINUX_HEADERS." " }
	    description "
This is the location of your RTAI and Linux kernel installation. It is normally
detected by the packages configure script and can be specified
with the argument --with-lxrt=path --with-linux=path  and modifyable in
the \"Detected Support Libraries->RTAI Installation\" 
package.
"
	}

#     cdl_option OROBLD_OS_LINUX_KERNEL {
# 	display "Target Linux Kernel Directory"
# 	description "
# Provide the location of the RTAI-patched linux kernel, for example, /usr/src/linux."
# 	flavor booldata
# 	default_value { "" }
# 	implements OROINT_OS_KERNEL_MODULE
#     }

    cdl_component OROSEM_OS_SCHEDTYPE {
	display "Scheduling Algorithm for Threads"
	description "
This option sets the default scheduling algorithm for the threads. 
See man sched_setscheduler for
more information on the available types. Set to SCHED_FIFO for
reliable applications ( functions not going in an endless loop), 
for non-realtime testing, set to SCHED_OTHER."
	flavor data
	default_value { "SCHED_OTHER" }
	legal_values { "SCHED_FIFO" "SCHED_RR" "SCHED_OTHER" }
    }

    cdl_component OROBLD_OS_ENABLE_LINUX_KERNEL {
	display "Build LXRT kernel Modules"
	description "
Enable this option when LXRT KERNEL MODULES need
to be build."
	parent CYGBLD_GLOBAL_OPTIONS
	flavor bool
	default_value 1
	implements OROINT_OS_KERNEL_MODULE

	cdl_option OROBLD_OS_LINUX_KERNEL {
	    display "Target Linux Kernel path"
	    flavor  data
	    no_define
 	    calculated { OROBLD_SUPPORT_RTAI_LINUX_KERNEL }
	    description "The path to the linux kernel when building kernel modules. For LXRT, this is set in 
	\"Detected Support Libraries->Kernel Directory\" package"
	}
    }


   cdl_component CYGBLD_GLOBAL_OPTIONS {
       display "Global build options"
       flavor none
       parent none
       description "
      Global build options including control over
      compiler flags, linker flags and choice of toolchain."

       cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
	   display "Global command prefix"
	   flavor  data
	   no_define
	   default_value { "" }
	   description "
        This option specifies the command prefix used when
        invoking the build tools."
       }

       cdl_option OROBLD_GLOBAL_CFLAGS_ADD {
	   display "User defined global compiler flags"
	   flavor  data
	   no_define
	   default_value {  "-pipe -Wall -Woverloaded-virtual" }
	   description   "
          This option allows you to override some global compiler flags.
The options you provide here will be appended to the CFLAGS variable below."
       }

       cdl_option CYGBLD_GLOBAL_LDFLAGS_ADD {
	   display "User defined linker flags"
	   flavor  data
	   no_define
	   default_value { "" }
	   description   "
          This option allows you to override the global linker flags.
          The options you provide here will be appended to the LDFLAGS variable.
          You can add additional library paths and flags here."
       }

       cdl_option OROBLD_OS_ARCHITECTURE {
	   display "Processor Target Architecture"
	   description "
This option will be added to the compiler flags.
Select here the processor architecture for which at least the
compiled code will run on."
	   flavor data
	   no_define
	   default_value { "pentium" }
	   legal_values { "pentium" "pentium2" "pentium3" "pentium4" "k6" "athlon" "athlon-xp" "athlon64" "none" }
       }

       cdl_option OROBLD_OS_PROCESSOR {
	   display "Tune to Processor Type"
	   description "
This option will be added to the compiler flags.
Select here the processor architecture at which the code will run
most tuned. We are forced to omit pentium/k6 processors, since this
would trigger non-thread-safe code generation when compiling. However,
your program will run on a pentium if selecting pentium4 or even athlon-xp for example."
	   flavor data
	   no_define
	   default_value { "pentium2" }
	   legal_values { "pentium2" "pentium3" "pentium4" "athlon" "athlon-xp" "athlon64" "none" }
       }

       cdl_option OROBLD_OS_ARCH {
	   display "Architecture Selection Macro"
	   description "
Depending on the above options (which modify compiler flags),
a different processor architecture is identified to enable processor
specific assembler instructions in Orocos."
	flavor data
	default_value { OROBLD_OS_ARCHITECTURE == "athlon64" ? "x86_64" : "i386" }
	legal_values { "x86_64" "i386" }
    }

    cdl_option CYGBLD_OS_CONFIG_SMP {
	    display "Build for SMP Systems"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor  bool
	    no_define
	    define CONFIG_SMP
	    default_value 0
	    description   "
Enable this flag if you want to use Orocos on SMP systems."
    }

    cdl_option CYGBLD_OS_COMPILER {
	    display "Compiler Features"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor  data
	    legal_values { "gcc2" "gcc3" "gcc4" }
	    default_value { OROPKG_SUPPORT_GCC_VERSION }
	    no_define
	    description   "
Here you can configure which compiler you use.
This may be detected automatically
in combination with the 'configure' script, providing
the option : CC=gcc-version"
    }

    cdl_component OROBLD_OS_OPTIMIZE {
	display "Optimization Strategy"
        description "
This option lets you control optimization of the overall Orocos
code. You can optimize for debugging or optimize for execution or compilation time. The difference
in application size and speed can be quite large when toggling this flag."
	flavor data
	    no_define
	default_value { "Execution" }
        legal_values { "Execution" "Debugging" "Compiling" }
	cdl_option OROBLD_OS_OPTIMIZE_DEBUGGING {
		display "Flags for debugging optimization"
        	description "
Compile with debugging info, no optimization flags and debug
code-checking on. Produces very large code size ( >100MB )."
		flavor data
		no_define
		active_if  { OROBLD_OS_OPTIMIZE == "Debugging" }
		default_value  { "-g -O0" }
	}
	cdl_option OROBLD_OS_OPTIMIZE_COMPILE {
		display "Flags for compile time optimization"
        	description "
Compile for fast compilation and allow debug macros.
Produces larger code size, but compiles very fast."
		flavor data
		no_define
		active_if { OROBLD_OS_OPTIMIZE == "Compiling" }
		default_value  { "-O" }
	}
	cdl_option OROBLD_OS_OPTIMIZE_EXECUTION {
		display "Flags for execution time optimization"
        	description "
Compile for fast execution and disable debugging macros.
This option delivers the smallest code size, but the longest
compilation times."
		flavor data
		no_define
		active_if { OROBLD_OS_OPTIMIZE == "Execution" }
		default_value  { "-O2 -DNDEBUG" }
	}
    }

	cdl_option CYGBLD_GLOBAL_CFLAGS {
	    display "Global compiler flags"
	    flavor  data
	    no_define
	    calculated { (OROBLD_OS_OPTIMIZE_EXECUTION ? OROBLD_OS_OPTIMIZE_EXECUTION : "").
		(OROBLD_OS_OPTIMIZE_DEBUGGING ? OROBLD_OS_OPTIMIZE_DEBUGGING : "").
		(OROBLD_OS_OPTIMIZE_COMPILE ? OROBLD_OS_OPTIMIZE_COMPILE : "").
		(OROBLD_OS_ARCHITECTURE == "none" ? "" :
		" -march=".OROBLD_OS_ARCHITECTURE).
		(OROBLD_OS_PROCESSOR == "none" ? "" : 
		(CYGBLD_OS_COMPILER == "gcc4" ? " -mtune=" : " -mcpu=" ).OROBLD_OS_PROCESSOR)." ".
		(OROBLD_OS_EXTRA_CFLAGS ? OROBLD_OS_EXTRA_CFLAGS : "")." ".
		"-D_REENTRANT ".
		(CYGBLD_OS_COMPILER == "gcc3" ? "" : "").
		(CYGBLD_OS_COMPILER == "gcc4" ? "-fvisibility-inlines-hidden " : "").
		OROBLD_GLOBAL_CFLAGS_ADD }
	    
	    description   "
This option controls the global compiler flags which
are used to compile all packages by
default. Individual packages may define
options which override these global flags. See also
the 'Optimization Strategy' to influence debugging or
execution speed compiler flags. 
You can not change these
flags but override them in the CYGBLD_GLOBAL_CFLAGS_ADD above.
Furthermore, depending on the compiler you selected, other flags may
be added."
	}

	cdl_option CYGBLD_GLOBAL_LDFLAGS {
	    display "Global linker flags"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor  data
	    no_define
	    default_value { "" }
	    description   "
This option controls the global linker flags. Individual
packages may define options which override these global flags."
	}

    cdl_option CYGBLD_LINKER_SCRIPT {
	display "Linker script"
	flavor data
	no_define
	calculated  { "" }
    }
    }

    cdl_option CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { "" }
    }

    cdl_option OROPKG_OS_LXRT_CFLAGS_REMOVE {
        display "Flags to remove for compiling"
        description "
RTAI/LXRT does not work well with -O3
"
        flavor data
        default_value { "-O3" }
    }

}
