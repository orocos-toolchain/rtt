
cdl_package OROPKG_DEVICE_DRIVERS_LOGICAL {
    display "C++ Interfaces to Logical Devices"
    parent OROPKG_DEVICE_DRIVERS

    include_dir device_drivers

    compile Axis.cxx DigitalInput.cxx DigitalOutput.cxx Drive.cxx DistanceSensor.cxx
    #compile SwitchEndLimit.cxx

}
