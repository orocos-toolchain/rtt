cdl_package OROPKG_KERNEL_COMPONENTS_PROCESS_CONTROL {
    parent OROPKG_KERNEL_COMPONENTS
    display "Signal and Process Control Components"
    description "
This package contains components for generating or
processing signals. It is usefull for rapid testing
hardware with one analog io card or generating/
controlling processes.
"
    requires OROPKG_CONTROL_KERNEL

    include_dir kernel_components

    compile SignalGenerator.cxx
    compile SignalTracker.cxx
    compile FeedForwardController.cxx
    compile P_Controller.cxx
    compile PID_Controller.cxx
}

