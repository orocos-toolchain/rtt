cdl_package OROPKG_DEVICE_DRIVERS_PORTS {
    display "Device Drivers for Standard IO Ports"
    description " This package contains a device
driver to access the parallel port.
"

    include_dir device_drivers
    include_files ParallelPort.hpp
    compile ParallelPort.cxx

    parent   OROPKG_DEVICE_DRIVERS
    requires OROPKG_DEVICE_DRIVERS
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
    requires OROINT_OS_LINUX_IOPERM

    cdl_component OROOPT_DEVICE_DRIVERS_PORTS_PARPORT_SCOPE {
	display "Use ParallelPort driver as Thread Scope"
	description "
When enabled, each Orocos thread will set a bit of this device
high or low to indicate its running status. The bit to thread
mapping is logged in the CoreLib Logger."
	flavor bool
	implements OROINT_DEVICE_INTERFACE_THREAD_SCOPE

	define_proc { 
	puts $::cdl_system_header "/***** proc output start *****/"
	puts $::cdl_system_header "#define ORODAT_DEVICE_DRIVERS_THREAD_SCOPE_INCLUDE <device_drivers/ParallelPort.hpp>"
	puts $::cdl_system_header "#define OROCLS_DEVICE_DRIVERS_THREAD_SCOPE_DRIVER ParallelPort"
	puts $::cdl_system_header "/****** proc output end ******/"
	}
    }

    cdl_option ORONUM_DEVICE_DRIVERS_PORTS_PARPORT {
	        display "Parallel Port Address"
		flavor data
        	default_value 0x378
    }

}