
cdl_package OROPKG_CORELIB_STATE {
    display "State infrastructure"
    description "
This package contains classes describing
States and how transitions between states
can be defined. It is used by the Execution
Package to form Machine States."

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    include_dir corelib

    compile StateInterface.cxx StateContext.cxx
}