    cdl_interface OROINT_DEVICE_DRIVERS_APCI2200 {
	flavor bool
    }

    cdl_option OROFUN_DEVICE_DRIVERS_APCI2200_LIB {
	no_define
	display "Calls to kernel module"
	description "
Only LXRT currently supports userspace code to call the kernel module." 
	calculated OROBLD_DEVICE_DRIVERS_APCI2200_KM && \
	    OROPKG_OS_LXRT
	implements OROINT_DEVICE_DRIVERS_APCI2200
	define_proc {
	    puts $::cdl_header "#define OROIMP_DEVICE_DRIVERS_APCI2200_T void"
	}
    }

cdl_option OROFUN_DEVICE_DRIVERS_APCI2200_IK {
    display "Built-in device driver"
    compile apci2200/apci2200.c
    calculated OROINT_OS_KERNEL
    implements OROINT_DEVICE_DRIVERS_APCI2200
	define_proc {
	    puts $::cdl_header "#define OROIMP_DEVICE_DRIVERS_APCI2200_T struct apci2200_device_t"
	}
}


    cdl_option OROBLD_DEVICE_DRIVERS_APCI2200_KM {
	display "Separate kernel module"
	description "
This option enables the build of a separate kernel module
when the target requires it."
	#requires !OROINT_OS_KERNEL
	calculated !OROINT_OS_KERNEL && OROINT_OS_KERNEL_MODULE
	make {
	    <PREFIX>/modules/apci2200.o: <PACKAGE>/src/apci2200/apci2200.c
	    $(CC) $(CFLAGS) -O2 -DMODULE -D__KERNEL__ -c $< -o $@
	}
    }
