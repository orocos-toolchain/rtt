cdl_package OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL_CARTESIAN {
    display "Control Kernel Components Cartesian Space Motion"
    description "
Components for 3D motion control, e.g. trajectory
planning and interpolation. An integrating simulator
is also provided for testing purposes.
"
    parent   OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL
    requires OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL
    requires OROPKG_GEOMETRY
    requires OROPKG_KINDYN

    include_dir control_kernel

    compile CartesianSensor.cxx
    compile CartesianEffector.cxx
    compile CartesianController.cxx
    compile CartesianGenerator.cxx
    compile CartesianEstimator.cxx
    compile CartesianPositionTracker.cxx
    compile CartesianProcess.cxx
}
