cdl_package OROPKG_DEVICE_DRIVERS_COMEDI {
    display "Comedi implementation of IO"

    cdl_option OROPKG_DEVICE_DRIVERS_COMEDI_CFLAGS_ADD {
        display "Comedi include path"
	description "The path is derived from the
detection of the packages configure script"
	flavor data
        default_value { "-I".OROBLD_SUPPORT_COMEDI_DIR }
    }

    include_dir comedi

    parent   OROPKG_DEVICE_DRIVERS

    requires OROPKG_SUPPORT_COMEDI
    requires OROPKG_DEVICE_DRIVERS
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
    requires OROPKG_DEVICE_INTERFACE_ENCODER
    
    compile ComediDevice.cxx ComediEncoder.cxx
}
