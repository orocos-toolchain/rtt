
cdl_package OROPKG_DEVICE_INTERFACE_LOGICAL {
    display "Device Interfaces Logical"

    description "
The Logical Device Interfaces represent Axis, Sensor etc
as logical devices instead of bare analog/digital IO."

    parent OROPKG_DEVICE_INTERFACE
    include_dir rtt/dev
    compile SensorInterface.cxx AxisInterface.cxx HomingInterface.cxx
}
