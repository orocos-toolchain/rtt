
cdl_package OROPKG_EXECUTION_PROGRAM_PROCESSOR {
    display "Program processing infrastructure"
    description "
A Package that provides realtime-safe program execution,
with each program statement represented by an object
which encapsulates the command to be executed."

    include_dir execution
    
    parent OROPKG_EXECUTION

    requires OROPKG_SUPPORT_BOOST_GRAPH
    requires OROPKG_SUPPORT_BOOST
    requires OROPKG_CORELIB_STATE

    compile StateContextBuilder.cxx
    compile VertexNode.cxx EdgeCondition.cxx ProgramGraph.cxx 
    compile CommandCounter.cxx  CommandIllegal.cxx  CommandString.cxx  
    compile ConditionBool.cxx  ConditionBoolDataSource.cxx  ConditionBoolProperty.cxx  ConditionComposite.cxx
    compile Processor.cxx
    compile AsynchCommandDecorator.cxx
    compile StateDescription.cxx
}
