cdl_package OROPKG_DEVICE_INTERFACE {
    display "C++ Hardware Device Interfaces"
}