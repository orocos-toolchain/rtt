
cdl_package OROPKG_CORELIB_PROPERTIES {
    display "Generic Property system"
    description "This package provides an implementation
       of any-type properties. Properties are
       an abstraction of the internal, configurable data of
       Components and can be read out and updated."

    include_dir corelib

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile PropertyBag.cxx  PropertySequence.cxx VectorComposition.cxx
    compile Property.cxx PropertyBase.cxx PropertyBagIntrospector.cxx
    compile OperationAcceptor.cxx

    cdl_option OROCLS_CORELIB_PROPERTIES_OPERATIONS {
	display "Property updating"
	description "Properties can be updated. Do not disable this option."
	active_if 1
	default_value 1
    }
}
