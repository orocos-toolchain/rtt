cdl_package OROPKG_GEOMETRY {
    display "Geometry library"
    description "
A Library representing the classes Vector, Rotation,
Frame, Twist, Wrench, Path, VelocityProfile, Trajectory
and others for 3D path planning, interpolation and kinematics"

    include_dir geometry
    
    compile debug_macros.cxx error_stack.cxx utility.cxx countingnumbers.cxx

    compile primitives/frame.cxx primitives/vector.cxx primitives/twist.cxx primitives/plane.cxx primitives/wrench.cxx
    compile primitives/rotation.cxx primitives/rframes.cxx primitives/rrframes.cxx primitives/rnframes.cxx
    compile primitives/plane.cxx

    compile primitives/path.cxx  primitives/path_circle.cxx  primitives/path_composite.cxx  primitives/path_cyclic_closed.cxx  
    compile primitives/path_line.cxx  primitives/path_point.cxx  primitives/path_roundedcomposite.cxx

    compile interpolation/velocityprofile.cxx
    compile interpolation/velocityprofile_dirac.cxx interpolation/velocityprofile_rect.cxx
    compile interpolation/velocityprofile_trap.cxx  interpolation/velocityprofile_traphalf.cxx
    compile interpolation/trajectory.cxx interpolation/trajectory_segment.cxx
    compile interpolation/rotational_interpolation.cxx  interpolation/rotational_interpolation_sa.cxx

    compile primitives/MotionProperties.cxx

#utility_newmat.cxx

    cdl_component OROPKG_GEOMETRY_3D {
	display "2D/3D Primitives Options"
	flavor none

	cdl_option OROSEM_GEOMETRY_ROTATION_PROPERTIES {
	    display "Rotation Property Format"
	    description "
Select this option to use Roll-Pitch-Yaw Angles when converting
Rotation Matrices to Properties or to use Euler Angles when converting
Rotation Matrices to Properties or to use
the lesser readable, but more accurate
Rotation Matrix (3x3 doubles) representation."
            flavor data
            default_value { "RPY" }
	    legal_values { "RPY" "EULER" "MATRIX" }
        }

	cdl_option OROPKG_GEOMETRY_3D_FRAMES_IO {
	    display "3D Primitives IO Marshalling"
	    description "
This enables the conversion of 3D primitives and trajectories to text streams
and back to binary format."
	    default_value 1
	    requires OROINT_OS_STDIOSTREAM
	    compile primitives/frames_io.cxx fileutils.cxx utility_io.cxx
	}

	cdl_option OROSEM_GEOMETRY_USE_EQUAL {
	    display "Use ORO_Geometry::Equal() for operator==()."
	    description "
Enable this option if you want the operator==() of frames, vectors,...
to use the Equal function, which compares the members of its arguments to a
'small' interval 'epsilon'. If disabled, the equality
operator for 'double' will be used on the members of these types"
            flavor bool
            default_value 1
        }

	cdl_option OROPKG_GEOMETRY_FRAMES_INLINE {
	    display "Try to inline small Frames methods."
	    description "
Enable this option if you want to inline small methods
for frame-related objects."
            flavor bool
            default_value 1
        }

    }
}

