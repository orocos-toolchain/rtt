
cdl_package OROPKG_EXECUTION_TASK_CONTEXT {
    display "Execution Task Context Infrastructure"
    description "
A Package that provides realtime-safe inter-task
communication and task browsing. A Task Context
contains the command-, method- and data-factories of that
task, a Processor which accepts commands and executes
task programs."

    include_dir execution
    
    parent OROPKG_EXECUTION

    requires OROPKG_EXECUTION
    requires OROPKG_EXECUTION_PROGRAM_PROCESSOR

    compile TaskContext.cxx
    compile AttributeRepository.cxx TaskAttribute.cxx 
    compile DataSourceFactoryInterface.cxx  GlobalDataSourceFactory.cxx
    compile GlobalCommandFactory.cxx
    compile CommandFactoryInterface.cxx
    compile PropertyLoader.cxx
    compile MapDataSourceFactory.cxx

}
