

cdl_package OROPKG_OS_LXRT {
    display "RTAI/LXRT OS Abstraction Layer"
    description "
Use this package if you want to compile 
Orocos for RTAI Realtime Userspace. It has
support for all packages used in Orocos."

    requires OROPKG_SUPPORT_RTAI

    include_dir os
    parent OROPKG_OS

    hardware

    compile PeriodicThread.cxx
    compile SingleThread.cxx
    compile MainThread.cxx
    compile main.cxx
    compile fosi.c

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB
    implements OROINT_OS_MAIN

    cdl_component OROCLS_OS_EVENT_INTERRUPT {
    }

    cdl_component OROSEM_OS_LXRT_SCHEDTYPE {
	display "Scheduling Algorithm for NOT realtime threads"
	description "
This option sets the scheduling algorithm for the threads
running in non-realtime. See man sched_setscheduler for
more information on the available types."
	flavor data
	default_value { "SCHED_OTHER" }
	legal_values { "SCHED_FIFO" "SCHED_RR" "SCHED_OTHER" }
    }

    cdl_option OROSEM_OS_LXRT_CHECK {
	display "Check LXRT calls for null pointers."
	description "
Enable to check for wrongly initialised pointers
when calling an LXRT function. You can disable this
for production code."
	flavor bool
	default_value 1
    }


    cdl_component CYGBLD_GLOBAL_OPTIONS {
	display "Global build options"
	flavor none
	parent CYGPKG_NONE
	description "
      Global build options including control over
      compiler flags, linker flags and choice of toolchain."

# 	cdl_option CYGBLD_GLOBAL_CFLAGS_ADD {
# 	    display "RTAI build directory include directive"
# 	    flavor data
# 	    default_value {"-I/usr/src/rtai"}
# 	    description "
# This is the location where rtai.h resides. It must
# point to a properly configured rtai installation."
# 	}
	cdl_option ORONUM_RTAI_VERSION {
	    display "RTAI version"
	    flavor data
	    #legal_values {"2" "3"}
	    calculated { OROBLD_SUPPORT_RTAI_VERSION }
	    description "
        Select the RTAI version you are using.
Legal values are 2 and 3. This value is detected by 
the packages configure script and modifyable in
the \"Detected Support Libraries->RTAI Installation\" 
package."
	}

	cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
	    display "Global command prefix"
	    flavor  data
	    no_define
	    default_value { "" }
	    description "
        This option specifies the command prefix used when
        invoking the build tools."
	}

	cdl_option CYGBLD_RTAIDIR {
	    display "RTAI directory"
	    flavor data
	    no_define
	    define -format="\\\"%s\/include\/config.h\\\"" ORO_RTAI_CONFIG
	    calculated { OROBLD_SUPPORT_RTAI_DIR }
	    description "
This is the location of your RTAI installation. It is normally
detected by the packages configure script and can be specified
with the argument --with-lxrt=path  and modifyable in
the \"Detected Support Libraries->RTAI Installation\" 
package.
"
	}

#     cdl_option OROBLD_OS_LINUX_KERNEL {
# 	display "Target Linux Kernel Directory"
# 	description "
# Provide the location of the RTAI-patched linux kernel, for example, /usr/src/linux."
# 	flavor booldata
# 	default_value { "" }
# 	implements OROINT_OS_KERNEL_MODULE
#     }

    cdl_component OROBLD_OS_ENABLE_LINUX_KERNEL {
	display "Build LXRT kernel Modules"
	description "
Enable this option when LXRT KERNEL MODULES need
to be build and set the correct path, for example
/usr/src/linux-rt"
	flavor bool
	default_value { 0 }
	implements OROINT_OS_KERNEL_MODULE

	cdl_option OROBLD_OS_LINUX_KERNEL {
	    display "Target Linux Kernel path"
	    flavor  data
	    no_define
	    default_value { "/usr/src/linux-rt" }
	    description "Provide the location of the RTAI-patched linux kernel, for example, /usr/src/linux-rt."
	}
    }
	cdl_option OROBLD_GLOBAL_CFLAGS_ADD {
	    display "User defined global compiler flags"
	    flavor  data
	    no_define
	    default_value { "" }
	    description   "
          This option allows you to override some global compiler flags.
The options you provide here will be appended to the CFLAGS variable.
You can add the '-g -O0' flags here for example."
	}

	cdl_option CYGBLD_GLOBAL_CFLAGS {
	    display "Global compiler flags"
	    flavor  data
	    no_define
	    calculated { " -pipe -Wall -Wnon-virtual-dtor -Woverloaded-virtual -O2 -I" . CYGBLD_RTAIDIR . "/include -march=". OROBLD_OS_ARCHITECTURE . " -mcpu=" .  OROBLD_OS_PROCESSOR . " " . OROBLD_GLOBAL_CFLAGS_ADD }
	    description   "
          This option shows the global compiler flags which
          are used to compile all packages by
          default. Individual packages may define
          options which override these global flags. You can not change these
          flags but override them in the CYGBLD_GLOBAL_CFLAGS_ADD"
	}

	cdl_option CYGBLD_GLOBAL_LDFLAGS_ADD {
	    display "User defined linker flags"
	    flavor  data
	    no_define
	    default_value { "" }
	    description   "
          This option allows you to override the global linker flags.
          The options you provide here will be appended to the LDFLAGS variable.
          You can add additional library paths and flags here."
	}

	cdl_option CYGBLD_GLOBAL_LDFLAGS {
	    display "Global linker flags"
	    flavor  data
	    no_define
	    calculated { " -L" . CYGBLD_RTAIDIR . "/lxrt/lib -L". CYGBLD_RTAIDIR. "/lib -llxrt" . CYGBLD_GLOBAL_LDFLAGS_ADD }
	    description   "
          This option controls the global linker flags. Individual
          packages may define options which override these global flags.
          You can not change these
          flags but override them in the CYGBLD_GLOBAL_LDFLAGS_ADD"
	}

    }

    cdl_option CYGBLD_LINKER_SCRIPT {
	display "Linker script"
	flavor data
	no_define
	calculated  { "" }
    }

    cdl_option CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { "" }
    }

}
