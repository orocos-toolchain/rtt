
cdl_package OROPKG_CORELIB_PROPERTIES_MARSHALLING {
    display "CoreLib Property Marshalling and Demarshalling"
    description "This package allows
to convert binary information to text (or another format) and vice
versa. There are marshallers for XML files, INI files and streaming
tables (for logging)."

    parent OROPKG_CORELIB_PROPERTIES
    requires OROPKG_CORELIB_PROPERTIES

    cdl_interface OROINT_CORELIB_PROPERTIES_MARSHALLING_FORMAT {
	requires { OROINT_CORELIB_PROPERTIES_MARSHALLING_FORMAT == 1 }
    }

    cdl_component OROPKG_CORELIB_PROPERTIES_MARSHALLING_DEFAULT {
	display "Defaul Marshalling Format"
	description "Select the default format which will be
used to read and write property files."
	
	flavor none
	no_define

	cdl_option OROPKG_CORELIB_PROPERTIES_MARSHALLING_CPF {
	    display "Component Property Format (XML) + Xerces"
	    description "
This Property format is standardised by the Object Management Group
(OMG) and is uses also in Corba 3 Components. It is quite readable
and powerful. It is very well tested within Orocos, but requires the heavy Xerses library."
	    requires OROPKG_SUPPORT_XERCESC
	    implements OROINT_CORELIB_PROPERTIES_MARSHALLING_FORMAT
	    default_value OROPKG_SUPPORT_XERCESC

	    define_proc { 
		puts $::cdl_header "/***** proc output start *****/"
		puts $::cdl_header "#define ORODAT_CORELIB_PROPERTIES_MARSHALLING_INCLUDE <rtt/marsh/CPFMarshaller.hpp>"
		puts $::cdl_header "#define OROCLS_CORELIB_PROPERTIES_MARSHALLING_DRIVER CPFMarshaller"
		puts $::cdl_header "#define ORODAT_CORELIB_PROPERTIES_DEMARSHALLING_INCLUDE <rtt/marsh/CPFDemarshaller.hpp>"
		puts $::cdl_header "#define OROCLS_CORELIB_PROPERTIES_DEMARSHALLING_DRIVER CPFDemarshaller"
		puts $::cdl_header "/****** proc output end ******/"
	    }

            compile CPFDemarshaller.cxx
	}

	cdl_option OROPKG_CORELIB_PROPERTIES_MARSHALLING_TINY_CPF {
	    display "Component Property Format (XML)"
	    description "
This Property format is standardised by the Object Management Group
(OMG) and is uses also in Corba 3 Components. It is quite readable
and powerful. It is very well tested within Orocos. This version uses
an internal 'TinyXML' library for minimal code size. It does not 
fully validate the correctness of the XML file (DTD)."
	    implements OROINT_CORELIB_PROPERTIES_MARSHALLING_FORMAT
	    default_value !OROPKG_SUPPORT_XERCESC

	    define_proc { 
		puts $::cdl_header "/***** proc output start *****/"
		puts $::cdl_header "#define ORODAT_CORELIB_PROPERTIES_MARSHALLING_INCLUDE <rtt/marsh/CPFMarshaller.hpp>"
		puts $::cdl_header "#define OROCLS_CORELIB_PROPERTIES_MARSHALLING_DRIVER CPFMarshaller"
		puts $::cdl_header "#define ORODAT_CORELIB_PROPERTIES_DEMARSHALLING_INCLUDE <rtt/marsh/TinyDemarshaller.hpp>"
		puts $::cdl_header "#define OROCLS_CORELIB_PROPERTIES_DEMARSHALLING_DRIVER TinyDemarshaller"
		puts $::cdl_header "/****** proc output end ******/"
	    }

            compile TinyDemarshaller.cxx
	    compile tinyxml.cxx tinyxmlparser.cxx tinyxmlerror.cxx tinystr.cxx
	}

    }
    include_dir rtt/marsh

    include_files CPFDemarshaller.hpp  INIMarshaller.hpp       Orocos1Demarshaller.hpp  SimpleDemarshaller.hpp  TableHeaderMarshaller.hpp  XMLDemarshaller.hpp  XMLRPCDemarshaller.hpp CPFDTD.hpp 
    include_files CPFMarshaller.hpp    MarshallerAdaptors.hpp  Orocos1Marshaller.hpp    SimpleMarshaller.hpp    TableMarshaller.hpp        XMLMarshaller.hpp    XMLRPCMarshaller.hpp
    include_files StreamProcessor.hpp EmptyHeaderMarshaller.hpp EmptyMarshaller.hpp 
    include_files TinyDemarshaller.hpp

    compile CPFDTD.cxx
}
