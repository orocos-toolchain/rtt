cdl_package OROPKG_OS_ECOS {
    display "OS Abstraction Layer eCos"
    description "
This package is used if you want to compile
Orocos for eCos, allowing hard
real-time userspace applications
"

    include_dir rtt/os
    parent OROPKG_OS

    compile fosi.c ecos_rec_mutex.c ecosthreads.cxx

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB

    define_proc {
        puts $::cdl_system_header "\#define CYGBLD_OS_TARGET_H   <pkgconf/os_ecos.h>"
    }

    cdl_option OROSEM_OS_ECOS_STACK_SIZE {
    display "Default stack size of ecos threads"
    description "
Set the stack size of the ecos threads
"
	flavor data
	# FIXME: For some f*cking reason, this doesn't work (although it
	# works with the net packages belonging to ecos 
	# default_value (CYGNUM_HAL_STACK_SIZE_TYPICAL*2)
	default_value 65536
    }

    # Fixme, inherit this from eCos
    cdl_component OROSEM_OS_SCHEDTYPE {
	display "Scheduling Algorithm for Threads"
	description "
This option sets the default scheduling algorithm for the threads.  
Only the CYGSEM_KERNEL_SCHED_MLQUEUE option is tested at this moment.
"
	flavor data
	default_value { "CYGSEM_KERNEL_SCHED_MLQUEUE" }
	legal_values { "CYGSEM_KERNEL_SCHED_MLQUEUE" "CYGSEM_KERNEL_SCHED_BITMAP" }
    }

    cdl_option ORONUM_OS_RTOS_HIGHEST_PRIORITY {
	display       "Highest possible priority"
	flavor data
	default_value    0
	description "All ecos schedulers use 0 as the highest
	priority, so you probably don't want to modify this variable"
    }

    cdl_option ORONUM_OS_RTOS_LOWEST_PRIORITY {
	display       "Lowest possible priority"
	flavor data
	default_value    CYGNUM_KERNEL_SCHED_PRIORITIES-1
	description "Lowest priority as configured by user. You
	probably don't want to modify this variable."
    }

    # Added by KG (reminder of kernel space modules?)
    # implements OROINT_OS_MAIN
    # requires OROPKG_SUPPORT_ECOS
}
