cdl_package OROPKG_KINDYN_ARCH {
    display "Kinematic and Dynamics Architectures"
    parent OROPKG_KINDYN
    requires OROPKG_KINDYN

    include_dir kindyn

    cdl_component OROPKG_KINDYN_ARCH_SERIAL321 {
	display "Serial 321 kinematics"
	description "Contains a number of kinematic
architectures for serial robots. The type of robot
is described in the Featherstone convention. Each letter denotes
the right-handed rotation around an axis of the robot base frame
of each respective joint. So Z***** means the first joint rotates
around the Z axis of the base frame. *X**** means the second joint
rotates around the X axis of the base frame, and so on."
	
	default_value 1

	compile serial321/ZXXDWH/SerialZXXDWH.cxx serial321/ZYYDWH/SerialZYYDWH.cxx
	compile serial321/ZXXDWH/ForJacZXXDWH.cxx  serial321/ZXXDWH/ForPosZXXDWH.cxx  serial321/ZXXDWH/ForVelZXXDWH.cxx  
	compile serial321/ZXXDWH/InvJacZXXDWH.cxx  serial321/ZXXDWH/InvPosZXXDWH.cxx  serial321/ZXXDWH/InvVelZXXDWH.cxx

    }
}

