cdl_package OROPKG_DEVICE_INTERFACE {
    display "Device Interfaces"
    description "
This package groups together all the hardware
abstraction interfaces. If you want to introduce
your hardware drivers into the Orocos framework,
they must be ported to these abstract C++ interfaces.

See the Device Drivers package for examples.
"
    include_files DeviceInterface.hpp
    include_dir rtt/dev

    cdl_interface OROINT_DEVICE_INTERFACE_THREAD_SCOPE {
	display "Support for a thread scope device driver"
	flavor data
	requires { OROINT_DEVICE_INTERFACE_THREAD_SCOPE <= 1 }
    }


}