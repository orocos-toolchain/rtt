
cdl_package OROPKG_CORELIB_PROPERTIES {
    display "Generic Property system"
    description "This package provides an implementation
       of a foreigntype-friendly properties. Properties are
       an abstraction of the internal, configurable data of
       components."

    include_dir corelib

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile PropertyBag.cxx  PropertySequence.cxx VectorComposition.cxx
    compile Property.cxx PropertyBase.cxx PropertyBagIntrospector.cxx

    cdl_option OROCLS_CORELIB_PROPERTIES_OPERATIONS {
	display "Cast-free property operations"
	description "This option enables the
           copy/mutate/update operations on the PropertyBase class."

	default_value 1
	compile OperationAcceptor.cxx
    }
}
