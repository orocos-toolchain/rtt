
cdl_package OROPKG_MATH {
    display "Math packages"
}