
cdl_package OROPKG_EXECUTION {
    display "Program logic execution Infrastructure"
}