
cdl_package OROPKG_CORELIB_CONDITIONS {
    display "CoreLib Condition abstraction interface definition"
    description "This package provides the ConditionInterface for
dynamic conditional execution of logic programs."

    include_dir corelib
    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile ConditionInterface.cxx
    compile ConditionDuration.cxx
    compile ConditionDSDuration.cxx
    compile ConditionOnce.cxx
    compile DataSourceCondition.cxx
}

