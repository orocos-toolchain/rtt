

cdl_package OROPKG_OS_GNULINUX {
    display "GNU/Linux OS abstraction layer"
    description "
This package is used if you want to compile
Orocos for 'User Space', not realtime. The
periodic threading support is very limited
and the package is mainly used for testing and
debugging other packages."

    include_dir os
    parent OROPKG_OS

    compile fosi.c
    compile ComponentThreaded.cxx
    compile SingleThread.cxx
    compile main.cxx

    implements OROINT_OS_STDCXXLIB
    implements OROINT_OS_KERNEL_MODULE

    cdl_component OROCLS_OS_EVENT_INTERRUPT {
	display "Interrupt driven event implementation (Dummy)"
	description "
This option causes an EventInterrupt class to be compiled,
but it will do nothing and will not react on interrupts."
	flavor bool
	implements OROINT_OS_EVENT_INTERRUPT
	compile EventInterrupt.cxx
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
	display "Global build options"
	flavor none
	parent CYGPKG_NONE
	description "
      Global build options including control over
      compiler flags, linker flags and choice of toolchain."

	cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
	    display "Global command prefix"
	    flavor  data
	    no_define
	    default_value { "" }
	    description "
        This option specifies the command prefix used when
        invoking the build tools."
	}

	cdl_option CYGBLD_GLOBAL_CFLAGS {
	    display "Global compiler flags"
	    flavor  data
	    no_define
	    default_value { "-g -pipe -Wall -Wstrict-prototypes -Woverloaded-virtual -Wnon-virtual-dtor -O2" }
	    description   "
          This option controls the global compiler flags which
          are used to compile all packages by
          default. Individual packages may define
          options which override these global flags."
	}

	cdl_option CYGBLD_GLOBAL_LDFLAGS {
	    display "Global linker flags"
	    flavor  data
	    no_define
	    default_value { "-g" }
	    description   "
          This option controls the global linker flags. Individual
          packages may define options which override these global flags."
	}
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
	display "Linker script"
	flavor data
	no_define
	calculated  { "" }
    }

    cdl_option CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { "" }
    }

}
