cdl_package OROPKG_OS {
    display "OS Abstraction Layer"
    description "
This Package groups operating system abstractions.
It defines a Thread, Mutex, IO and the capabilities
of the system for which Orocos is compiled. You
can only select one OS Package which is called the
'target'."

    include_dir os
    
    compile startstop.cxx
    compile StartStopManager.cxx
    compile Mutex.cxx

    cdl_option OROBLD_OS_AGNOSTIC {
	display "Hide system includes from Orocos headers."
	description "
When enabled, Orocos OS headers will not expose non standard system file
includes to the library user. In other words, every OS function call is
wrapped and they are not inlined. This makes it easier to compile
applications with Orocos headers, since no extra include paths must be
added (like /usr/realtime). Also Built-in assembly instructions
will be used instead of the system header files.
"
	flavor bool
        default_value 1
    }

    cdl_option OROCLS_OS_MINIMAL_STREAMS {
	display "Minimal streams implementation"
	description "
This provides an <iostream> like implementation of
streams, but suitable for hard realtime at the cost
of generality (so it is less configurable as the 
std C++ library). It resides in the rt_std namespace."
	flavor bool
	default_value 1
	compile rtstreams.cxx
	compile rtconversions.cxx  rtctype.cxx
    }

    cdl_option OROFUN_OS_ALTERNATE_RTTI {
	display "Alternate C++ Run Time Type Info (EXP)"
	description "
Enable to compile a C++ RTTI implementation, based on the
gcc compilers implementation. Only use if your target's
C++ libraries have no RTTI support *and* use with care."
	flavor bool
	default_value 0
	compile rt_tinfo.cxx rt_tinfo2.cxx
	active_if OROCFG_CORELIB_EXPERIMENTAL
    }

    cdl_option OROBLD_OS_ARCHITECTURE {
	display "Processor Target Architecture"
        description "
This option will be added to the compiler flags.
Select here the processor architecture for which at least the
compiled code will run on."
	flavor data
	default_value { "pentium" }
        legal_values { "pentium" "pentium2" "pentium3" "pentium4" "k6" "athlon" "athlon-xp" }
    }

    cdl_option OROBLD_OS_PROCESSOR {
	display "Tune to Processor Type"
        description "
This option will be added to the compiler flags.
Select here the processor architecture at which the code will run
most tuned. We are forced to omit pentium/k6 processors, since this
would trigger non-thread-safe code generation when compiling. However,
your program will run on a pentium if selecting pentium4 or even athlon-xp for example."
	flavor data
	default_value { "pentium2" }
        legal_values { "pentium2" "pentium3" "pentium4" "athlon" "athlon-xp" }
    }

    # we need exactly one OS_TARGET
    cdl_interface OROINT_OS_TARGET {
	display "Target Operating System"
	flavor bool
	requires OROINT_OS_TARGET == 1
    }

    cdl_interface OROINT_OS_GLOBAL_CRT {
	display "Target calls global constructors"
	flavor bool
	requires OROINT_OS_GLOBAL_CRT <= 1
	define HAVE_MANUAL_CRT
    }

    cdl_interface OROINT_OS_MAIN {
	display "Target which simulates a main function"
	flavor bool
	requires OROINT_OS_MAIN <= 1
	define HAVE_MANUAL_MAIN
    }

    cdl_interface OROINT_OS_EVENT_INTERRUPT {
	display "Support for interrupt based Events"
	flavor bool
    }

    cdl_interface OROINT_OS_STDCXXLIB {
	display "Support for the Standard C++ Library"
	flavor bool
	implements OROINT_OS_STDVECTOR
	implements OROINT_OS_STDLIST
	implements OROINT_OS_STDMAP
	implements OROINT_OS_STDSTRING
	implements OROINT_OS_STDIOSTREAM
    }

    cdl_interface OROINT_OS_STDVECTOR {
	display "Vector of the Standard C++ Library"
	flavor bool
    }

    cdl_interface OROINT_OS_STDLIST {
	display "List of the Standard C++ Library"
	flavor bool
    }

    cdl_interface OROINT_OS_STDQUEUE {
	display "Queue of the Standard C++ Library"
	flavor bool
    }

    cdl_interface OROINT_OS_STDMAP {
	display "Map of the Standard C++ Library"
	flavor bool
    }

    cdl_interface OROINT_OS_STDSTRING {
	display "String of the Standard C++ Library"
	flavor bool
    }

    cdl_interface OROINT_OS_STDIOSTREAM {
	display "IOStreams of the Standard C++ Library"
	flavor bool
    }

    cdl_interface OROINT_OS_KERNEL {
	display "Inside-kernel interface"
	flavor bool
    }

    cdl_interface OROINT_OS_KERNEL_MODULE {
	display "Kernel module loader support"
	flavor bool
    }

    cdl_interface OROINT_OS_RECURSIVE_MUTEX {
	display "Support for recursive mutex"
	flavor bool
    }
}
