cdl_package OROPKG_GEOMETRY {
    display "Geometry library"
    description "
A Library representing the classes Vector, Rotation,
Frame, Twist, Wrench, Path, VelocityProfile, Trajectory
and others for 3D path planning and interpolation."

    include_dir geometry
    
    compile debug_macros.cxx error_stack.cxx utility.cxx countingnumbers.cxx

#utility_newmat.cxx

    cdl_component OROPKG_GEOMETRY_3D {
	display "3D Primitives"
	default_value 1

	cdl_option OROPKG_GEOMETRY_3D_FRAMES {
	    display "3D Frames, Twists, Wrenches"
	    description "
This contains implementations of 3D Vector, Rotation, Frame,
Twist and Wrench"
	    default_value 1
	    compile primitives/frame.cxx primitives/vector.cxx primitives/twist.cxx primitives/plane.cxx primitives/wrench.cxx
	    compile primitives/rotation.cxx primitives/rframes.cxx primitives/rrframes.cxx primitives/rnframes.cxx
	    compile primitives/plane.cxx
	}

	cdl_option OROSEM_GEOMETRY_EULERPROPERTIES {
	    display "Use Euler ZYX Angles for Properties"
	    description "
Enable this option to use Euler Angles when converting
Rotation Matrices to Properties or vice versa. When
disabled, The lesser readable, but more accurate
Rotation Matrix (3x3) will be marshalled."
            flavor bool
            default_value 1
            active_if OROPKG_GEOMETRY_3D_FRAMES
        }

	cdl_option OROPKG_GEOMETRY_3D_FRAMES_IO {
	    display "3D IO conversions"
	    description "
This enables the conversion of 3D primitives to text streams
and back to binary format."
	    default_value 1
	    requires OROINT_OS_STDIOSTREAM
	    compile primitives/frames_io.cxx fileutils.cxx utility_io.cxx
	}

	cdl_option OROPKG_GEOMETRY_3D_PROPERTIES {
	    display "Geometry Property Support"
	    description "
This enables the conversion of 3D primitives within Properties
to basic Properties and back. You will need this if you want to
use Property<Frame> and the like as a property."
	    default_value 1
	    requires OROINT_OS_STDIOSTREAM
	    compile primitives/MotionProperties.cxx
	}

    }

    cdl_component OROPKG_GEOMETRY_PRIMITIVES {
	display "Path Primitives"
	description "
This includes Path_Line, Path_Point, Path_Circle,
Path_Cyclic_Closed, Path_Composite and Path_RoundedComposite"
	default_value 1
	active_if OROPKG_GEOMETRY_3D_FRAMES
	compile primitives/path.cxx  primitives/path_circle.cxx  primitives/path_composite.cxx  primitives/path_cyclic_closed.cxx  
	compile primitives/path_line.cxx  primitives/path_point.cxx  primitives/path_roundedcomposite.cxx
    }

    cdl_component OROPKG_GEOMETRY_INTERPOLATION {
	display "Interpolation algorithms"
	description "
Velocity profile planning and trajectory composition"
	flavor bool
	default_value 1
	active_if OROPKG_GEOMETRY_3D_FRAMES && OROPKG_GEOMETRY_PRIMITIVES

	compile interpolation/velocityprofile.cxx
        compile interpolation/velocityprofile_dirac.cxx interpolation/velocityprofile_rect.cxx
        compile interpolation/velocityprofile_trap.cxx  interpolation/velocityprofile_traphalf.cxx
	compile interpolation/trajectory.cxx  interpolation/trajectory_composite.cxx  interpolation/trajectory_segment.cxx
	compile interpolation/rotational_interpolation.cxx  interpolation/rotational_interpolation_sa.cxx

    }
}

