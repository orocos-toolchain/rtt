cdl_package OROPKG_CONTROL_KERNEL_COMPONENTS {
    display "Control Kernel components"
    description "
Components for Control Kernels. This parent
package contains some common, application
independent Components like a console command reader
and a console output component."

    parent   OROPKG_CONTROL_FRAMEWORK
    requires OROPKG_CONTROL_FRAMEWORK
    requires OROPKG_CONTROL_KERNEL
    requires OROPKG_SUPPORT_READLINE

    include_dir control_kernel

    compile HMIConsoleOutput.cxx HMIConsoleInput.cxx
    compile HMIReadline.cxx
}
