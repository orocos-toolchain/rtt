cdl_package OROPKG_DEVICE_DRIVERS_CANOPEN {
    display "Device Drivers CANOpen implementation based on CANPie"
    description "
This package was made for controlling a Beckhoff
based CANOpen bus for an industrial partner."

    include_dir can

    parent   OROPKG_DEVICE_DRIVERS

    requires OROPKG_DEVICE_DRIVERS
    requires OROPKG_DEVICE_DRIVERS_CANPIE
    requires OROINT_DEVICE_DRIVERS_CP_CORE
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
    requires OROPKG_DEVICE_INTERFACE_ENCODER
    
    compile CAN.cxx
    compile CANPieController.cxx
    compile BeckhoffCANCoupler.cxx
}