
cdl_package OROPKG_CORELIB_ACTIVITIES {
    display "CoreLib Periodic Activity/Thread Infrastructure"
    description "
This packages allows you to create Periodic Activities and (realtime) Threads.
Activities of equal priority are serialised in the same thread.
Therefore, Orocos specifies in advance three types of threads
with different priorities and semantics. Each thread has a different
type of periodic activity associated with it. 
"
    include_dir rtt

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile PeriodicActivity.cxx
    compile TimerThread.cxx
    compile SimulationThread.cxx SimulationActivity.cxx NonPeriodicActivity.cxx
    compile TimerSequencer.cxx TimerOneShot.cxx TimerLockFree.cxx
    compile CoreRunnableInterface.cxx SlaveActivity.cxx
}

