
cdl_package OROPKG_EXECUTION_PROGRAM_PARSER {
    display "Execution Script-to-Program parser"
    description "
Converts text files (scripts) to realtime binary programs
for the Program Processor using the Boost::Spirit
library. It takes a lot of time to compile, but
is very powerful."

    include_dir execution

    parent OROPKG_EXECUTION

    compile Types.cxx Operators.cxx
    compile CommonParser.cxx
    compile parse_exception.cxx
    compile StateGraphParser.cxx
    compile ArgumentsParser.cxx ConditionParser.cxx ExpressionParser.cxx Parser.cxx
    compile ValueParser.cxx CommandParser.cxx ProgramGraphParser.cxx ValueChangeParser.cxx
    compile DataSourceCondition.cxx DataSourceCommand.cxx 
    compile ParsedStateMachine.cxx
    compile StateMachineBuilder.cxx
    compile PeerParser.cxx 
    compile PropertyParser.cxx 
    compile FunctionFactory.cxx
    compile TaskBrowser.cxx
    compile ProgramLoader.cxx
    compile GenericTaskContext.cxx
    compile StatementProcessor.cxx

    requires OROPKG_SUPPORT_BOOST
    requires OROPKG_SUPPORT_BOOST_GRAPH 
    requires OROPKG_SUPPORT_BOOST_PARSER
    requires OROPKG_SUPPORT_READLINE
    requires OROPKG_CORELIB_PROPERTIES
    requires OROPKG_EXECUTION
    requires OROPKG_EXECUTION_PROGRAM_PROCESSOR
    requires OROPKG_EXECUTION_TASK_CONTEXT

    cdl_option OROPKG_EXECUTION_PROGRAM_PARSER_CFLAGS_REMOVE {
        display "Flags to remove for compiling"
        description "
Normally we compile without debugging info because
it generates huge object files.
"
        flavor data
        default_value { "-g" }
    }
}
