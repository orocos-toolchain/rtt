
cdl_package OROPKG_DEVICE_DRIVERS_LOGICAL {
    display "Device Drivers C++ Interfaces to Logical Devices"
    description "
This package has some 'common' implementations
for addressing single channels of devices. For
example, a DigitalInput channel, an Axis or
an AnalogDrive. They interface with Device Interface
classes."
    parent OROPKG_DEVICE_DRIVERS
    requires OROPKG_CORELIB_EVENTS

    include_dir rtt/dev

    compile Axis.cxx SimulationAxis.cxx DigitalInput.cxx DigitalOutput.cxx AnalogDrive.cxx AbsoluteEncoderSensor.cxx IncrementalEncoderSensor.cxx
}
