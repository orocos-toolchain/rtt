
cdl_package OROPKG_EXECUTION_TASK_CONTEXT {
    display "Execution Task Context Infrastructure"
    description "
A Package that provides realtime-safe inter-task
communication and task browsing. A Task Context
contains the command-, method- and data-factories of that
task, a Processor which accepts commands and executes
task programs."

    include_dir rtt
    
    parent OROPKG_EXECUTION

    requires OROPKG_EXECUTION
    requires OROPKG_CORELIB
    requires OROPKG_CORELIB_PROPERTIES
    requires OROPKG_CORELIB_COMMANDS

    cdl_component OROPKG_EXECUTION_ENGINE {
	display "Execution Engine Configuration"
	description "Enable or disable various parts
of the standard ExecutionEngine"
	flavor none
	cdl_component OROPKG_EXECUTION_ENGINE_EVENTS {
	    display "Enable Event Processor"
	    description "If disabled, the EventProcessor is removed from the ExecutionEngine."
	    default_value OROPKG_CORELIB_EVENTS
	    active_if OROPKG_CORELIB_EVENTS
	    flavor bool
	    compile EventService.cxx
	    compile EventC.cxx
            compile ConnectionC.cxx
	}
	cdl_component OROPKG_EXECUTION_ENGINE_COMMANDS {
	    display "Enable Command Processor"
	    description "If disabled, the CommandProcessor is removed from the ExecutionEngine."
	    default_value 1
	    active_if OROPKG_EXECUTION_PROGRAM_PROCESSOR
	    flavor bool
	}
	cdl_component OROPKG_EXECUTION_ENGINE_PROGRAMS {
	    display "Enable Program Processor"
	    description "If disabled, the ProgramProcessor is removed from the ExecutionEngine."
	    default_value 1
	    flavor bool
	}
	cdl_component OROPKG_EXECUTION_ENGINE_STATEMACHINES {
	    display "Enable StateMachine Processor"
	    description "If disabled, the StateMachineProcessor is removed from the ExecutionEngine."
	    default_value 1
	    active_if OROPKG_EXECUTION_PROGRAM_PROCESSOR
	    flavor bool
	}

    }

    compile TaskContext.cxx
    compile AttributeRepository.cxx
    compile PropertyLoader.cxx
    compile ExecutionEngine.cxx
    compile CommandC.cxx
    compile MethodC.cxx
    compile ScriptingAccess.cxx
    compile TryCommand.cxx
    compile ConnectionInterface.cxx
    compile PortInterface.cxx
    compile TaskCore.cxx
}
