
cdl_package OROPKG_CORELIB_EVENTS {
    display "CoreLib Synchronous-Asynchronous Event system"
    description "
This package provides an Event implementation for
synchronous and asynchronous event handling."

    include_dir rtt
    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    implements OROINT_CORELIB_EVENT_INTERFACE
    implements OROINT_CORELIB_COMPLETION_INTERFACE

    compile EventProcessor.cxx
    compile signal_base.cxx
    compile Handle.cxx
    compile CompletionProcessor.cxx

}