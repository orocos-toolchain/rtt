
cdl_package OROPKG_CORELIB_REPORTING {
    display "CoreLib Reporting and Logging Infrastructure"
    description "This package adds binary to text reporting
of internal data in a separate thread. It is mainly used for
logging and data gathering. See the README for a short 
description of the nomenclature. Also, contains the Orocos
Logger implementation for tracking system configuration."

    include_dir corelib

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile ReportWriter.cxx
    compile ReportCollectorInterface.cxx PropertyExporter.cxx
    compile Logger.cxx

    requires OROPKG_CORELIB_PROPERTIES

    cdl_component OROBLD_CORELIB_REPORTING_LOGGING {
	display "Configure Logging Messages"
	no_define
	flavor none
	cdl_option OROBLD_CORELIB_REPORTING_DISABLE_LOGGING {
	    display "Disable all Logging."
	    define OROBLD_DISABLE_LOGGING
	    description "
Enable this option to disable the Logger. No logging messages
will be displayed or written to the orocos.log file."
	    flavor bool
	    default_value 0
	}

	cdl_option OROBLD_CORELIB_REPORTING_PRINTF_LOGGING {
	    display "Log using printf/fprintf"
	    define OROSEM_PRINTF_LOGGING
	    active_if !OROBLD_CORELIB_REPORTING_DISABLE_LOGGING
	    description "
Enable this option to use only printf / fprintf for logging instead of
iostream and fstream (std::cout, ...)"
	    flavor bool
	    default_value 0
	}

	cdl_option OROBLD_CORELIB_REPORTING_FILE_LOGGING {
	    display "Log to orocos.log"
	    define OROSEM_FILE_LOGGING
	    active_if !OROBLD_CORELIB_REPORTING_DISABLE_LOGGING
	    description "
Enable this option to write the logs to a file, orocos.log, as well."
	    flavor bool
	    default_value 1
	}

	cdl_option OROBLD_CORELIB_REPORTING_REMOTE_LOGGING {
	    display "Store logs in memory for retrieval."
	    define OROSEM_REMOTE_LOGGING
	    active_if !OROBLD_CORELIB_REPORTING_DISABLE_LOGGING
	    description "
Enable this option to store the logs IN MEMORY for later retrieval
by a different (remote) component. Does not use printf nor iostreams."
	    flavor bool
	    default_value 1
	}

	cdl_option ORONUM_CORELIB_REPORTING_LOGGING_BUFFER {
	    display "Maximum log lines held in memory."
	    define ORONUM_LOGGING_BUFSIZE
	    active_if !OROBLD_CORELIB_REPORTING_DISABLE_LOGGING && OROBLD_CORELIB_REPORTING_REMOTE_LOGGING
	    description "
When remote logging is enabled, the log messages are stored in
memory until fetched by a client. In order to avoid memory
exhaustion, a maximum number of messages is stored. If this
number is exceeded, a FIFO principle is used to remove the
oldest messages."
	    flavor data
	    default_value 1000
	}
    }

}
