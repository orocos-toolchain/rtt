cdl_package OROPKG_KERNEL_COMPONENTS {
    display "Control Kernel components"
    description "
Components for Control Kernels. This parent
package contains some common, application
independent Components."

    requires OROPKG_CONTROL_KERNEL

    include_dir kernel_components

    compile HMIConsoleOutput.cxx HMIConsoleInput.cxx
    compile HMIReadline.cxx
}
