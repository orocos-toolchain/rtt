

cdl_package OROPKG_OS_LXRT {
    display "OS Abstraction Layer RTAI/LXRT"
    description "
Use this package if you want to compile 
Orocos for RTAI Realtime Userspace. It has
support for all packages used in Orocos."

    requires OROPKG_SUPPORT_RTAI

    include_dir os
    parent OROPKG_OS

    hardware

    compile MainThread.cxx
    compile fosi.c

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB
    implements OROINT_OS_MAIN
    implements OROINT_OS_LINUX_IOPERM

    cdl_option OROSEM_OS_LXRT_CHECK {
	display "Check LXRT calls for null pointers."
	description "
Enable to check for wrongly initialised pointers
when calling an LXRT function. You can disable this
for production code."
	flavor bool
	default_value 1
    }

    cdl_option OROSEM_OS_LXRT_PERIODIC {
	display "Run RTAI Scheduler in periodic mode"
	description "
Enable to use the periodic mode of the RTAI scheduler
instead of the 'one-shot' scheduler. You need to provide
the periodic scheduler execution period in seconds (s). Leave this
disabled if unsure."
	flavor booldata
	default_value 0
	define ORODAT_OS_LXRT_PERIODIC_TICK
    }


	cdl_option ORONUM_RTAI_VERSION {
	    display "RTAI version"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor data
	    #legal_values {"2" "3"}
	    calculated { OROBLD_SUPPORT_RTAI_VERSION }
	    description "
        Select the RTAI version you are using.
Legal values are 2 and 3. This value is detected by 
the packages configure script and modifyable in
the \"Detected Support Libraries->RTAI Installation\" 
package."
	}

	cdl_option CYGBLD_RTAIDIR {
	    display "RTAI directory"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor data
	    no_define
	    define -format="\\\"%s\/include\/config.h\\\"" ORO_RTAI_CONFIG
	    calculated { OROBLD_SUPPORT_RTAI_DIR }
	    description "
This is the location of your RTAI installation. It is normally
detected by the packages configure script and can be specified
with the argument --with-lxrt=path  and modifyable in
the \"Detected Support Libraries->RTAI Installation\" 
package.
"
	}

#     cdl_option OROBLD_OS_LINUX_KERNEL {
# 	display "Target Linux Kernel Directory"
# 	description "
# Provide the location of the RTAI-patched linux kernel, for example, /usr/src/linux."
# 	flavor booldata
# 	default_value { "" }
# 	implements OROINT_OS_KERNEL_MODULE
#     }

    cdl_component OROBLD_OS_ENABLE_LINUX_KERNEL {
	display "Build LXRT kernel Modules"
	description "
Enable this option when LXRT KERNEL MODULES need
to be build and set the correct path, for example
/usr/src/linux-rt"
	parent CYGBLD_GLOBAL_OPTIONS
	flavor bool
	default_value { 0 }
	implements OROINT_OS_KERNEL_MODULE

	cdl_option OROBLD_OS_LINUX_KERNEL {
	    display "Target Linux Kernel path"
	    flavor  data
	    no_define
	    default_value { "/usr/src/linux-rt" }
	    description "Provide the location of the RTAI-patched linux kernel, for example, /usr/src/linux-rt."
	}
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
	display "Linker script"
	flavor data
	no_define
	calculated  { "" }
    }

    cdl_option CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { "" }
    }

}
