
cdl_package OROPKG_CORELIB_EVENTS {
    display "CoreLib Synchronous-Asynchronous Event system"
    description "
This package provides an Event implementation for
synchronous and asynchronous event handling."

    include_dir corelib
    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    implements OROINT_CORELIB_EVENT_INTERFACE

    compile EventProcessor.cxx
    compile signal_base.cxx
    compile Handle.cxx

    cdl_option OROSEM_CORELIB_EVENTS_ASYN {
	display "Enable asynchronous event completion."
	description "
This means a part of the event (called the completion)
can be deferred to another thread."
	flavor bool
	compile CompletionProcessor.cxx
	implements OROINT_CORELIB_COMPLETION_INTERFACE
    }

    cdl_option OROSEM_CORELIB_EVENTS_AUTOSTART {
	display "Automatically start the CompletionProcessor"
	description "
This option will enable starting the CompletionProcessor thread
automatically in the background so that the application does
no longer have to do so."
	flavor bool
	default_value 1
    }

    cdl_component OROPKG_CORELIB_EVENTS_CP {
	display "Completion Processor Properties"
	description "
The Completion Processor is a thread which processes
periodically deferred completion requests of events."
	flavor none
	requires OROSEM_CORELIB_EVENTS_ASYN
	
	cdl_option ORODAT_CORELIB_EVENTS_CP_NAME {
	    display "The name of the completion processor"
	    description "
The name must be unique with respect to other threads."
	    flavor data
	    default_value {"\"CompletionProcessor\""}
	    #legal_values string
	}
	cdl_option ORONUM_CORELIB_EVENTS_CP_PERIOD {
	    display "The periodicity of the completion processor in seconds"
	    description "
Indicates the time between processing two completion requests.
Since the request is inherently deferred (delayed), this value should mostly not
be smaller then 0.01 second."
	    flavor data
	    default_value 0.05
	    #legal_values positive number
	}
	cdl_option ORONUM_CORELIB_EVENTS_CP_PRIORITY {
	    display "The priority of the completion processor"
            description "
Every thread needs a priority. The completion processor is by
default not realtime though, so this value is less important."
	    flavor data
	    default_value 5
	    #legal_values positive number
	}
    }
}