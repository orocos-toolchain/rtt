
cdl_package OROPKG_DEVICE_INTERFACE_IO {
    display "Device Interfaces to A/D IO cards"
    description "
The interfaces are for Digital Input cards,
Digital Output cards, Analog Input cards and
Analog Output cards."

    parent OROPKG_DEVICE_INTERFACE

    include_dir rtt/dev

    compile io.cxx
}