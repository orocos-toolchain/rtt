
cdl_interface OROINT_DEVICE_DRIVERS_APCI1032 {
	flavor bool
    }


cdl_option OROFUN_DEVICE_DRIVERS_APCI1032_LIB {
    no_define
    display "Calls to kernel module"
    description "
Only LXRT currently supports userspace code to call the kernel module." 
    calculated OROBLD_DEVICE_DRIVERS_APCI1032_KM && \
	OROPKG_OS_LXRT
    implements OROINT_DEVICE_DRIVERS_APCI1032
    define_proc {
	puts $::cdl_header "#define OROIMP_DEVICE_DRIVERS_APCI1032_T void"
    }
}

cdl_option OROFUN_DEVICE_DRIVERS_APCI1032_IK {
    display "Built-in device driver"
    compile apci1032/apci1032.c
    calculated OROINT_OS_KERNEL
    implements OROINT_DEVICE_DRIVERS_APCI1032
    define_proc {
	puts $::cdl_header "#define OROIMP_DEVICE_DRIVERS_APCI1032_T struct apci1032_device_t"
    }
}


cdl_option OROBLD_DEVICE_DRIVERS_APCI1032_KM {
    display "Separate kernel module"
    description "
This option enables the build of a separate kernel module
when the target requires it."
    #requires !OROINT_OS_KERNEL
    calculated !OROINT_OS_KERNEL && OROINT_OS_KERNEL_MODULE
    make {
	<PREFIX>/modules/apci1032.o: <PACKAGE>/src/apci1032/apci1032.c
	$(CC) $(CFLAGS) -O2 -DMODULE -D__KERNEL__ -c $< -o $@
    }
}

cdl_option OROCLS_DEVICE_DRIVERS_APCI1032_EVENTS {
    display "Event based input change notification"
    flavor bool
    requires OROCFG_CORELIB_EXPERIMENTAL && OROINT_CORELIB_EVENT_INTERFACE
    description "
Enable to make the SwitchDigitalInapci1032 a Preemptible Task
which will fire an event if the inputs change."
}
