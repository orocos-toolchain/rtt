
cdl_package OROPKG_EXECUTION_PROGRAM_PARSER {
    display "Script-to-Program parser"
    description "
Converts text files (scripts) to realtime binary programs
for the Program Processor using the Boost::Spirit
library. It takes a lot of time to compile, but
is very powerful."

    include_dir execution

    parent OROPKG_EXECUTION

    compile CommonParser.cxx
    compile parse_exception.cxx
    compile StateGraphParser.cxx
    compile ArgumentsParser.cxx ConditionParser.cxx ExpressionParser.cxx Parser.cxx
    compile ValueParser.cxx CommandParser.cxx ProgramGraphParser.cxx ValueChangeParser.cxx
    compile Types.cxx DataSourceCondition.cxx Operators.cxx CommandFactoryInterface.cxx
    compile GlobalCommandFactory.cxx DataSource.cxx DataSourceFactoryInterface.cxx 
    compile GlobalDataSourceFactory.cxx
    compile ParsedStateContext.cxx
    compile PeerParser.cxx
    compile ParsedValue.cxx ValueRepository.cxx

    requires OROPKG_SUPPORT_BOOST
    requires OROPKG_SUPPORT_BOOST_GRAPH 
    requires OROPKG_EXECUTION_PROGRAM_PROCESSOR

    cdl_option OROPKG_EXECUTION_PROGRAM_PARSER_CFLAGS_REMOVE {
        display "Flags to remove for compiling"
        description "
Normally we compile without debugging info because
it generates huge object files.
"
        flavor data
        default_value { "-g" }
    }
}
