cdl_package OROPKG_KERNEL_COMPONENTS_MOTION_CONTROL_AXIS {
    display "Multi Axis control components"
    description "
Components for 1D Axis motion control, e.g. trajectory
planning and interpolation.
"
    parent OROPKG_KERNEL_COMPONENTS_MOTION_CONTROL
    requires OROPKG_KERNEL_COMPONENTS_MOTION_CONTROL

    requires OROPKG_CONTROL_KERNEL
    requires OROPKG_GEOMETRY
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
    requires OROPKG_DEVICE_INTERFACE_LOGICAL

    include_dir kernel_components

    compile AxisSensor.cxx AxisEffector.cxx
    compile AxisPositionGenerator.cxx
}
