cdl_package OROPKG_KERNEL_COMPONENTS_MOTION_CONTROL {
    display "Motion Control Components"
    description "
Components for 1D or 3D motion control.
"
    parent OROPKG_KERNEL_COMPONENTS
    requires OROPKG_KERNEL_COMPONENTS

    requires OROPKG_CONTROL_KERNEL
}
