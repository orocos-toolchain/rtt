cdl_package OROPKG_KERNEL_COMPONENTS_MOTION_CONTROL {
    display "Motion control components"
    description "
Components for 1D or 3D motion control, e.g. trajectory
planning and interpolation, axis-level control,...
A special Sensor, Generator and Effector are included
for multi-Axis motion control.
"
    parent OROPKG_KERNEL_COMPONENTS

    requires OROPKG_CONTROL_KERNEL

    include_dir kernel_components

    compile sensor/AxisSensor.cxx effector/AxisEffector.cxx

    compile sensor/CartesianNSSensor.cxx
    compile effector/CartesianNSEffector.cxx
    compile controller/CartesianNSController.cxx
    compile generator/CartesianNSGenerator.cxx
    compile estimator/CartesianNSEstimator.cxx

    compile generator/AxisPositionGenerator.cxx generator/CartesianPositionTracker.cxx
}
