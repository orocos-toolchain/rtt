cdl_package OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL_AXIS {
    display "Control Kernel Components Motion Control Multi Axis"
    description "
Components for 1D Axis motion control, e.g. trajectory
planning and interpolation.
"
    parent   OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL
    requires OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL
    requires OROPKG_GEOMETRY
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
    requires OROPKG_DEVICE_INTERFACE_LOGICAL

    include_dir control_kernel

    compile AxisSensor.cxx AxisEffector.cxx
    compile AxisPositionGenerator.cxx
}
