cdl_package OROPKG_DEVICE_DRIVERS_COMEDI {
    display "Device Drivers Comedi implementation of IO"

    cdl_option OROPKG_DEVICE_DRIVERS_COMEDI_CFLAGS_ADD {
        display "Comedi include path"
	description "The path is derived from the
detection of the packages configure script"
	flavor data
        default_value { "-I".OROBLD_SUPPORT_COMEDI_DIR }
    }

    include_dir rtt/dev

    parent   OROPKG_DEVICE_DRIVERS

    requires OROPKG_SUPPORT_COMEDI
    requires OROPKG_DEVICE_DRIVERS
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
    requires OROPKG_DEVICE_INTERFACE_ENCODER
    
    compile ComediDevice.cxx ComediEncoder.cxx
    compile ComediSubDeviceDOut.cxx ComediSubDeviceAOut.cxx
    compile ComediSubDeviceDIn.cxx ComediSubDeviceAIn.cxx

    cdl_component OROOPT_DEVICE_DRIVERS_COMEDI_THREAD_SCOPE {
	display "Use Comedi driver as Thread Scope"
	description "
When enabled, each Orocos thread will set a bit of this device
high or low to indicate its running status. The bit to thread
mapping is logged in the CoreLib Logger."
	flavor bool
	implements OROINT_DEVICE_INTERFACE_THREAD_SCOPE

	cdl_option ORODAT_DEVICE_DRIVERS_COMEDI_THREAD_SCOPE_MINOR {
	        display "Thread Scope Comedi device minor"
		description "
The minor device number which you want to use for the scope.
To use /dev/comedi0 , enter 0."
		flavor data
        	default_value 0
	}

	cdl_option ORODAT_DEVICE_DRIVERS_COMEDI_THREAD_SCOPE_SUBDEVICE {
	        display "Thread Scope Comedi subdevice"
		description "
The comedi subdevice which you want to use for the scope. It
must be a digital output subdevice."
		flavor data
        	default_value 0
	}

	define_proc { 
	puts $::cdl_system_header "/***** proc output start *****/"
	puts $::cdl_system_header "#define ORODAT_DEVICE_DRIVERS_THREAD_SCOPE_INCLUDE <rtt/dev/ComediThreadScope.hpp>"
	puts $::cdl_system_header "#define OROCLS_DEVICE_DRIVERS_THREAD_SCOPE_DRIVER ComediThreadScope"
	puts $::cdl_system_header "/****** proc output end ******/"
	}
    }

}
