
cdl_package OROPKG_CORELIB_TIMING {
    display "CoreLib Time measurement infrastructure"
    description "This package contains the 
TimeService which will be used to keep track of system
time and defines time conversions."

    include_dir rtt

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile TimeService.cxx
}
