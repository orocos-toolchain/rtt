
cdl_package OROPKG_CORELIB_BUFFERS {
    display "CoreLib Communication buffers"
    description "
This package contains the lock-free communication buffers
for local (in-process) data exchange. A lock-free single
linked list and pointer queue is provided as well."

    include_dir rtt
    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile BufferLockFree.cxx
    compile ListLockFree.cxx
    compile DataObjectInterfaces.cxx	
}