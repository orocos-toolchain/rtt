
cdl_package OROPKG_CORELIB_PROPERTIES {
    display "CoreLib Generic Property system"
    description "This package provides an implementation
       of any-type properties. Properties are
       an abstraction of the internal, configurable data of
       Components and can be read out and updated."

    include_dir rtt

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB
    requires OROPKG_CORELIB_COMMANDS

    compile PropertyBag.cxx  PropertySequence.cxx VectorComposition.cxx
    compile Property.cxx PropertyBase.cxx PropertyBagIntrospector.cxx

}
