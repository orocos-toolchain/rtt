cdl_package OROPKG_CONTROL_KERNEL_COMPONENTS_HARDWARE {
    display "Control Kernel Components Hardware access"
    description "
Easy to use Components that can use device drivers
which implement the Orocos Device Interface. The 
Components will read or write to kernel DataObjects
and provide commands for the Program Execution Extension.
The package contains a Sensor and an Effector
Component."

    parent   OROPKG_CONTROL_KERNEL_COMPONENTS
    requires OROPKG_CONTROL_KERNEL_COMPONENTS

    include_dir control_kernel

    compile GenericSensor.cxx GenericEffector.cxx

    requires OROPKG_CONTROL_KERNEL
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
}
