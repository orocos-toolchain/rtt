cdl_package OROPKG_SIGNAL_PROCESSING {
    display "Signal Processing Library"
    description "
A Library for generating or modifying analog or digital signals.
It is only for demonstrative purposes now and needs to be filled
in by a non Orocos project. It just contains a sine generator."

    include_dir signal_processing
}

