
cdl_package OROPKG_EXECUTION {
    display "Program logic execution Infrastructure"
    description "
This Package groups infrastructure for parsing and
executing realtime program logic in the Orocos Framework."
}