

cdl_package OROPKG_OS_XENOMAI {
    display "OS Abstraction Layer Xenomai 2.0"
    description "
This package is used if you want to compile
Orocos for Xenomai 2.0, allowing
real-time userspace applications"

    include_dir os
    parent OROPKG_OS

    compile fosi.c

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB
    implements OROINT_OS_LINUX_IOPERM

    requires OROPKG_SUPPORT_XENOMAI

    hardware

    cdl_component OROBLD_OS_ENABLE_LINUX_KERNEL {
	display "Build Linux kernel Modules"
	description "
Enable this option when Linux KERNEL MODULES need
to be build and set the correct path, for example
/usr/src/linux"
	parent CYGBLD_GLOBAL_OPTIONS
	flavor bool
	default_value 1
	implements OROINT_OS_KERNEL_MODULE

	cdl_option OROBLD_OS_LINUX_KERNEL {
	    display "Target Linux Kernel path"
	    flavor  data
	    no_define
	    default_value { OROBLD_SUPPORT_FUSION_LINUX_KERNEL }
	    description "The target linux path."
	}
    }

	cdl_option OROBLD_OS_EXTRA_CFLAGS {
	    display "Fusion Include Directory"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor data
	    no_define
	    calculated { "-I".OROBLD_SUPPORT_FUSION_DIR."/include -I".OROBLD_SUPPORT_FUSION_LINUX_HEADERS." " }
	    description "
This is the location of your Xenomai and Linux kernel installation. It is normally
detected by the packages configure script and can be specified
with the argument --with-xenomai=path --with-linux=path  and modifyable in
the \"Detected Support Libraries->Xenomai Installation\" 
package.
"
	}

    cdl_option CYGBLD_LINKER_SCRIPT {
	display "Linker script"
	flavor data
	no_define
	calculated  { "" }
    }

    cdl_option CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { "" }
    }

}
