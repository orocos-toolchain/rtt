

cdl_package OROPKG_OS_GNULINUX {
    display "OS Abstraction Layer GNU/Linux"
    description "
This package is used if you want to compile
Orocos for 'User Space', not realtime. The
periodic threading support is very limited
and the package is mainly used for testing and
debugging other packages."

    include_dir os
    parent OROPKG_OS

    compile fosi.c

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB
    implements OROINT_OS_LINUX_IOPERM


    cdl_component OROBLD_OS_ENABLE_LINUX_KERNEL {
	display "Build Linux kernel Modules"
	description "
Enable this option when Linux KERNEL MODULES need
to be build and set the correct path, for example
/usr/src/linux"
	parent CYGBLD_GLOBAL_OPTIONS
	flavor bool
	default_value 1
	implements OROINT_OS_KERNEL_MODULE

	cdl_option OROBLD_OS_LINUX_KERNEL {
	    display "Target Linux Kernel path"
	    flavor  data
	    no_define
	    default_value { "********SET LINUX KERNEL PATH IN GLOBAL BUILD OPTIONS OR DISABLE 'Build Linux Kernel Modules'********" }
	    description "The target linux path."
	}
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
	display "Linker script"
	flavor data
	no_define
	calculated  { "" }
    }

    cdl_option CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { "" }
    }

}
