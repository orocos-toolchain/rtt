cdl_package OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL_N_AXIS { 
    display "Control Kernel Components Motion Control N-Axis"
    description "
Components for N-Axis motion control, e.g. trajectory
planning and interpolation.
"
    parent   OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL
    requires OROPKG_CONTROL_KERNEL_COMPONENTS_MOTION_CONTROL
    requires OROPKG_GEOMETRY
    requires OROPKG_KINDYN
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO
    requires OROPKG_DEVICE_INTERFACE_LOGICAL

    include_dir control_kernel

    compile nAxesControllerPos.cxx nAxesControllerPosVel.cxx nAxesControllerVel.cxx
    compile nAxesControllerCartesianPosVel.cxx nAxesControllerCartesianPos.cxx nAxesControllerCartesianVel.cxx
    compile nAxesEffectorVel.cxx nAxesEffectorCartesianVel.cxx
    compile nAxesGeneratorPos.cxx nAxesGeneratorSin.cxx nAxesGeneratorCartesianPos.cxx nAxesGeneratorVel.cxx nAxesGeneratorCartesianSin.cxx
    compile nAxesSensorPos.cxx nAxesSensorCartesianPos.cxx nAxesSensorCartesianPosForce.cxx  nAxesSensorForcesensor.cxx 
}
