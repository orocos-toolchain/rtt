
cdl_package OROPKG_CORELIB_COMMANDS {
    display "CoreLib Command abstraction interface definition"
    description "
      This Package is required for logical program execution.
      It provides utilities and the interface for the CommandInterface."

    include_dir rtt

    parent OROPKG_CORELIB
    requires OROPKG_CORELIB

    compile CommandNOP.cxx
    compile DataSourceCommand.cxx

}
