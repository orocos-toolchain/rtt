
cdl_package OROPKG_EXECUTION_PROGRAM_PARSER {
    display "Script-to-Program parser"
    include_dir execution

    parent OROPKG_EXECUTION

    compile ArgumentsParser.cxx ConditionParser.cxx ExpressionParser.cxx Parser.cxx
    compile ValueParser.cxx CommandParser.cxx ProgramParser.cxx ValueChangeParser.cxx
    compile Types.cxx DataSourceCondition.cxx Operators.cxx CommandFactoryInterface.cxx

    requires OROPKG_SUPPORT_BOOST
}