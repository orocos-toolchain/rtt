

cdl_package OROPKG_OS_XENOMAI {
    display "OS Abstraction Layer Xenomai 2.0"
    description "
This package is used if you want to compile
Orocos for Xenomai 2.0, allowing
real-time userspace applications"

    include_dir os
    parent OROPKG_OS

    compile fosi.c
    compile MainThread.cxx

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB
    implements OROINT_OS_MAIN
    implements OROINT_OS_LINUX_IOPERM

    requires OROPKG_SUPPORT_XENOMAI

    hardware

    cdl_component OROBLD_OS_ENABLE_LINUX_KERNEL {
	display "Build Linux kernel Modules"
	description "
Enable this option when Linux KERNEL MODULES need
to be build and set the correct path, for example
/usr/src/linux"
	parent CYGBLD_GLOBAL_OPTIONS
	flavor bool
	default_value 1
	implements OROINT_OS_KERNEL_MODULE

	cdl_option OROBLD_OS_LINUX_KERNEL {
	    display "Target Linux Kernel path"
	    flavor  data
	    no_define
	    default_value { OROBLD_SUPPORT_XENOMAI_LINUX_KERNEL }
	    description "The target linux path."
	}
    }

    cdl_option OROSEM_OS_XENO_CHECK {
	display "Check Xenomai calls for null pointers."
	description "
Enable to check for wrongly initialised pointers
when calling an Xenamai function. You can disable this
for production code."
	flavor bool
	default_value 1
    }

    cdl_option OROSEM_OS_XENO_PERIODIC {
	display "Run Xenomai Scheduler in periodic mode"
	description "
Enable to use the periodic mode of the Xenomai scheduler
instead of the 'one-shot' scheduler. You need to provide
the periodic scheduler execution period in seconds (s). Leave this
disabled if unsure."
	flavor booldata
	default_value 0
	define ORODAT_OS_XENO_PERIODIC_TICK
    }

	cdl_option OROBLD_OS_EXTRA_CFLAGS {
	    display "Xenomai Include Directory"
	    parent CYGBLD_GLOBAL_OPTIONS
	    flavor data
	    no_define
	    calculated { "-I".OROBLD_SUPPORT_XENOMAI_DIR."/include -I".OROBLD_SUPPORT_XENOMAI_LINUX_HEADERS." " }
	    description "
This is the location of your Xenomai and Linux kernel installation. It is normally
detected by the packages configure script and can be specified
with the argument --with-xenomai=path --with-linux=path  and modifyable in
the \"Detected Support Libraries->Xenomai Installation\" 
package.
"
	}

    cdl_option CYGBLD_LINKER_SCRIPT {
	display "Linker script"
	flavor data
	no_define
	calculated  { "" }
    }

    cdl_option CYGHWR_MEMORY_LAYOUT {
	display "Memory layout"
	flavor data
	no_define
	calculated { "" }
    }

}
