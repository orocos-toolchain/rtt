cdl_package OROPKG_CONTROL_KERNEL_COMPONENTS_KINEMATICS {
    display "Control Kernel Components for Kinematics"
    description "
Kinematic Components for Control Kernels. This
package contains process components for doing kinematic
calculations and kinematic state stracking."

    parent   OROPKG_CONTROL_KERNEL_COMPONENTS
    requires OROPKG_CONTROL_KERNEL_COMPONENTS
    requires OROPKG_CONTROL_KERNEL

    include_dir control_kernel

    include_files KinematicProcess.hpp
    compile KinematicProcess.cxx
}
