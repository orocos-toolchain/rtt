cdl_package OROPKG_KERNEL_COMPONENTS_PROCESS_CONTROL {
    parent OROPKG_KERNEL_COMPONENTS
    display "Signal and Process Control Components"
    description "
This package contains components for generating or
processing signals. It is usefull for rapid testing
hardware with one analog io card or generating/
controlling processes. It contains P, PID and
FeedForward Controllers. Multi Channel signals
can be generated using the signal Generator
and a signal tracker Generator Components.
Works very good in conjunction with the Motion Control
and Hardware Components.
"
    requires OROPKG_KERNEL_COMPONENTS

    include_dir kernel_components

    compile SignalGenerator.cxx
    compile SignalTracker.cxx
    compile FeedForwardController.cxx
    compile P_Controller.cxx
    compile PID_Controller.cxx
}

