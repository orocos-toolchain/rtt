cdl_package OROPKG_CONTROL_KERNEL_SERVER {
    display "Control Kernel CORBA Server"
    description "
A CORBA server which allows your kernel to be used with the KernelClient GUI.
"
    parent   OROPKG_CONTROL_FRAMEWORK
    requires OROPKG_CONTROL_FRAMEWORK

    include_dir control_kernel

    make_object {
	src/kernelserver.o : $(REPOSITORY)/$(PACKAGE)/src/KernelInterface.idl
	tao_idl $(REPOSITORY)/$(PACKAGE)/src/KernelInterface.idl -o src
	touch $@
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/src/kernelserver.cxx -o src/$(OBJECT_PREFIX)_kernelserver.o
    }

    make_object {
	src/KernelInterfaceI.o : $(REPOSITORY)/$(PACKAGE)/src/KernelInterface.idl
	touch $@
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/src/KernelInterfaceI.cxx -o src/$(OBJECT_PREFIX)_KernelInterfaceI.o
    }

    make_object {
	src/KernelInterfaceS.o : $(REPOSITORY)/$(PACKAGE)/src/KernelInterface.idl
	touch $@
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c src/KernelInterfaceS.cpp -o src/$(OBJECT_PREFIX)_KernelInterfaceS.o
    }

    make_object {
	src/KernelInterfaceS_T.o : $(REPOSITORY)/$(PACKAGE)/src/KernelInterface.idl
	touch $@
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c src/KernelInterfaceS_T.cpp -o src/$(OBJECT_PREFIX)_KernelInterfaceS_T.o
    }

    make_object {
	src/KernelInterfaceC.o : $(REPOSITORY)/$(PACKAGE)/src/KernelInterface.idl
	touch $@
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c src/KernelInterfaceC.cpp -o src/$(OBJECT_PREFIX)_KernelInterfaceC.o
    }

#    compile KernelInterfaceI.cxx
#    compile kernelserver.cxx
    compile directkernelinterface.cxx
    compile kernelinterface.cxx

}
