cdl_package OROPKG_KERNEL_COMPONENTS {
    display "Control Kernel components"
    description "
Components for Control Kernels. This parent
package contains some common, application
independent Components like a console command reader
and a console output component."

    requires OROPKG_CONTROL_KERNEL

    include_dir kernel_components

    compile HMIConsoleOutput.cxx HMIConsoleInput.cxx
    compile HMIReadline.cxx
}
