cdl_package OROPKG_CORBA {
    display "Control Task CORBA Framework"
    description "
This package allows to tranparantly setup remote Tasks
and connect to them from local tasks. Only minor CORBA/RPC
knowledge is required to use this framework.
"
    requires OROPKG_EXECUTION_TASK_CONTEXT
    requires OROPKG_SUPPORT_CORBA

    implements OROINT_OS_CORBA

    cdl_option OROPKG_CORBA_CFLAGS_ADD {
        display "ACE/TAO include path"
	description "The path is derived from the
detection of the packages configure script"
	flavor data
        default_value { "-I".OROBLD_SUPPORT_ACE_DIR." -I".OROBLD_SUPPORT_TAO_DIR." -I".OROBLD_SUPPORT_TAO_DIR."/orbsvcs" }
    }

    include_dir rtt/corba
    include_files ApplicationServer.hpp
    include_files ControlTaskProxy.hpp ControlTaskServer.hpp ExpressionProxy.hpp  ScriptingAccessProxy.hpp
    include_files ExpressionServer.hpp CORBAExpression.hpp ActionProxy.hpp CommandProxy.hpp
    include_files Operations.idl OperationsC.h OperationsS.h OperationsC.inl OperationsS.inl OperationsS_T.h OperationsS_T.inl OperationsS_T.cpp OperationsI.h
    include_files ControlTask.idl ControlTaskC.h ControlTaskS.h ControlTaskC.inl ControlTaskS.inl ControlTaskS_T.h ControlTaskS_T.inl ControlTaskS_T.cpp ControlTaskI.h
    include_files OperationInterface.idl OperationInterfaceC.h OperationInterfaceS.h OperationInterfaceC.inl OperationInterfaceS.inl OperationInterfaceS_T.h OperationInterfaceS_T.inl OperationInterfaceS_T.cpp OperationInterfaceI.h
    include_files CosPropertyServiceI.h
    include_files CorbaMethodFactory.hpp CorbaCommandFactory.hpp CorbaConversion.hpp 
    include_files OrocosTypesC.h OrocosTypesC.inl GeometryConversion.hpp
    include_files GeometryC.h GeometryC.inl
    include_files Attributes.idl AttributesC.h AttributesS.h AttributesC.inl AttributesS.inl AttributesS_T.h AttributesS_T.inl AttributesS_T.cpp AttributesI.h
    include_files ScriptingAccess.idl ScriptingAccessC.h ScriptingAccessS.h ScriptingAccessC.inl ScriptingAccessS.inl ScriptingAccessS_T.h ScriptingAccessS_T.inl ScriptingAccessS_T.cpp ScriptingAccessI.h
    include_files Corba.hpp CorbaPort.hpp Services.hpp 
    include_files CorbaDataObject.hpp CorbaDataObjectProxy.hpp
    include_files CorbaBuffer.hpp CorbaBufferProxy.hpp POAUtility.h
    include_files DataFlow.idl DataFlowC.h DataFlowS.h DataFlowC.inl DataFlowS.inl DataFlowS_T.h DataFlowS_T.inl DataFlowS_T.cpp DataFlowI.h
    include_files Services.idl ServicesC.h ServicesS.h ServicesC.inl ServicesS.inl ServicesS_T.h ServicesS_T.inl ServicesS_T.cpp ServicesI.h


#     make_object {
# 	src/kernelserver.o : $(REPOSITORY)/$(PACKAGE)/ControlTask.idl $(REPOSITORY)/$(PACKAGE)/src/kernelserver.cxx
# 	tao_idl $(REPOSITORY)/$(PACKAGE)/src/KernelInterface.idl -o src
# 	touch $@
# 	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/src/kernelserver.cxx -o src/$(OBJECT_PREFIX)_kernelserver.o
#     }

    cdl_option OROPKG_CORBA_GEOMETRY {
	display "Geometry Corba Support"
	description "When the geometry package is used,
            Corba support will be enabled for the Frame, Vector, Twist,... types."
	flavor bool
	calculated OROPKG_GEOMETRY

	make_object {
	    GeometryC.o : $(REPOSITORY)/$(PACKAGE)/include/Geometry.idl
	    $(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/include/GeometryC.cpp -o $(OBJECT_PREFIX)_GeometryC.o
	    touch $@
	}
    }

    make_object {
	OrocosTypesC.o : $(REPOSITORY)/$(PACKAGE)/OrocosTypes.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/OrocosTypesC.cpp -o $(OBJECT_PREFIX)_OrocosTypesC.o
	touch $@
    }

    make_object {
	src/ControlTaskI.o : $(REPOSITORY)/$(PACKAGE)/ControlTask.idl $(REPOSITORY)/$(PACKAGE)/src/ControlTaskI.cpp
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/src/ControlTaskI.cpp -o src/$(OBJECT_PREFIX)_ControlTaskI.o
	touch $@
    }

    make_object {
	ControlTaskS.o : $(REPOSITORY)/$(PACKAGE)/ControlTask.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/ControlTaskS.cpp -o $(OBJECT_PREFIX)_ControlTaskS.o
	touch $@
    }

    make_object {
	ControlTaskC.o : $(REPOSITORY)/$(PACKAGE)/ControlTask.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/ControlTaskC.cpp -o $(OBJECT_PREFIX)_ControlTaskC.o
	touch $@
    }

    #AttributeInterface
    make_object {
	src/AttributesI.o : $(REPOSITORY)/$(PACKAGE)/Attributes.idl $(REPOSITORY)/$(PACKAGE)/src/AttributesI.cpp
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/src/AttributesI.cpp -o src/$(OBJECT_PREFIX)_AttributesI.o
	touch $@
    }

    make_object {
	AttributesS.o : $(REPOSITORY)/$(PACKAGE)/Attributes.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/AttributesS.cpp -o $(OBJECT_PREFIX)_AttributesS.o
	touch $@
    }

    make_object {
	AttributesC.o : $(REPOSITORY)/$(PACKAGE)/Attributes.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/AttributesC.cpp -o $(OBJECT_PREFIX)_AttributesC.o
	touch $@
    }

	#Operations Servers
    make_object {
	src/OperationsI.o : $(REPOSITORY)/$(PACKAGE)/Operations.idl $(REPOSITORY)/$(PACKAGE)/src/OperationsI.cpp
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/src/OperationsI.cpp -o src/$(OBJECT_PREFIX)_OperationsI.o
	touch $@
    }

    make_object {
	OperationsS.o : $(REPOSITORY)/$(PACKAGE)/Operations.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/OperationsS.cpp -o $(OBJECT_PREFIX)_OperationsS.o
	touch $@
    }

    make_object {
	OperationsC.o : $(REPOSITORY)/$(PACKAGE)/Operations.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/OperationsC.cpp -o $(OBJECT_PREFIX)_OperationsC.o
	touch $@
    }

    # OperationInterface servers
    make_object {
	src/OperationInterfaceI.o : $(REPOSITORY)/$(PACKAGE)/OperationInterface.idl $(REPOSITORY)/$(PACKAGE)/src/OperationInterfaceI.cpp
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/src/OperationInterfaceI.cpp -o src/$(OBJECT_PREFIX)_OperationInterfaceI.o
	touch $@
    }

    make_object {
	OperationInterfaceS.o : $(REPOSITORY)/$(PACKAGE)/OperationInterface.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/OperationInterfaceS.cpp -o $(OBJECT_PREFIX)_OperationInterfaceS.o
	touch $@
    }

    make_object {
	OperationInterfaceC.o : $(REPOSITORY)/$(PACKAGE)/OperationInterface.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/OperationInterfaceC.cpp -o $(OBJECT_PREFIX)_OperationInterfaceC.o
	touch $@
    }

    #ScriptingAccess
    make_object {
	src/ScriptingAccessI.o : $(REPOSITORY)/$(PACKAGE)/ScriptingAccess.idl $(REPOSITORY)/$(PACKAGE)/src/ScriptingAccessI.cpp
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/src/ScriptingAccessI.cpp -o src/$(OBJECT_PREFIX)_ScriptingAccessI.o
	touch $@
    }

    make_object {
	ScriptingAccessS.o : $(REPOSITORY)/$(PACKAGE)/ScriptingAccess.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/ScriptingAccessS.cpp -o $(OBJECT_PREFIX)_ScriptingAccessS.o
	touch $@
    }

    make_object {
	ScriptingAccessC.o : $(REPOSITORY)/$(PACKAGE)/ScriptingAccess.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/ScriptingAccessC.cpp -o $(OBJECT_PREFIX)_ScriptingAccessC.o
	touch $@    }

    #DataFlow
    make_object {
	src/DataFlowI.o : $(REPOSITORY)/$(PACKAGE)/DataFlow.idl $(REPOSITORY)/$(PACKAGE)/src/DataFlowI.cpp
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/src/DataFlowI.cpp -o src/$(OBJECT_PREFIX)_DataFlowI.o
	touch $@
    }

    make_object {
	DataFlowS.o : $(REPOSITORY)/$(PACKAGE)/DataFlow.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/DataFlowS.cpp -o $(OBJECT_PREFIX)_DataFlowS.o
	touch $@
    }

    make_object {
	DataFlowC.o : $(REPOSITORY)/$(PACKAGE)/DataFlow.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/DataFlowC.cpp -o $(OBJECT_PREFIX)_DataFlowC.o
	touch $@    }

    #Services
    make_object {
	ServicesS.o : $(REPOSITORY)/$(PACKAGE)/Services.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/ServicesS.cpp -o $(OBJECT_PREFIX)_ServicesS.o
	touch $@
    }

    make_object {
	ServicesC.o : $(REPOSITORY)/$(PACKAGE)/Services.idl
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -Isrc/ -O2 -c $(REPOSITORY)/$(PACKAGE)/ServicesC.cpp -o $(OBJECT_PREFIX)_ServicesC.o
	touch $@    }


    #CosPropertyService
    make_object {
	src/CosPropertyServiceI.o : $(REPOSITORY)/$(PACKAGE)/src/CosPropertyServiceI.cpp
	$(CC) $(CFLAGS) $(INCLUDE_PATH) -O2 -c $(REPOSITORY)/$(PACKAGE)/src/CosPropertyServiceI.cpp -o src/$(OBJECT_PREFIX)_CosPropertyServiceI.o
	touch $@
    }


    compile ApplicationServer.cxx
    compile ControlTaskProxy.cxx
    compile ControlTaskServer.cxx
    compile ExpressionProxy.cxx
    compile ExpressionServer.cxx
    compile ActionProxy.cxx
    compile CommandProxy.cxx
    compile CorbaConversion.cxx
    compile ScriptingAccessProxy.cxx
    compile CorbaDataObject.cxx CorbaDataObjectProxy.cxx
    compile CorbaBuffer.cxx CorbaBufferProxy.cxx
    compile Services.cxx POAUtility.cxx
}
