
cdl_package OROPKG_EXECUTION_PROGRAM_PROCESSOR {
    display "Program processing infrastructure"
    include_dir execution
    
    parent OROPKG_EXECUTION

    requires OROPKG_CORELIB_STATE

    compile VertexNode.cxx EdgeCondition.cxx ProgramGraph.cxx 
    compile CommandCounter.cxx  CommandIllegal.cxx  CommandString.cxx  
    compile ConditionBool.cxx  ConditionBoolDataSource.cxx  ConditionBoolProperty.cxx  ConditionComposite.cxx
    compile Processor.cxx  ProcessorState.cxx  ProcessorStateConfig.cxx  ProcessorStateExec.cxx  ProcessorStateInit.cxx  ProcessorStateLoad.cxx  
    compile Rule.cxx  RulesAbortList.cxx  RulesCheckList.cxx  RulesList.cxx
    compile SystemContext.cxx  SystemState.cxx
    compile AsynchCommandDecorator.cxx
}