cdl_package OROPKG_CONTROL_KERNEL_COMPONENTS_PROCESS_CONTROL {
    display "Control Kernel Components for Signal and Process Control"
    description "
This package contains components for generating or
processing signals. It is usefull for rapid testing
hardware with one analog io card or generating/
controlling processes. It contains P, PID and
FeedForward Controllers. Multi Channel signals
can be generated using the signal Generator
and a signal tracker Generator Components.
Works very good in conjunction with the Motion Control
and Hardware Components.
"
    parent   OROPKG_CONTROL_KERNEL_COMPONENTS
    requires OROPKG_CONTROL_KERNEL_COMPONENTS

    include_dir control_kernel

    compile SignalGenerator.cxx
    compile SignalTracker.cxx
    compile FeedForwardController.cxx
    compile P_Controller.cxx
    compile PID_Controller.cxx
}

