
cdl_package OROPKG_EXECUTION_PROGRAM_PROCESSOR {
    display "Execution Program processing infrastructure"
    description "
A Package that provides realtime-safe program execution,
with each program statement represented by an object
which encapsulates the command to be executed."

    include_dir execution
    
    parent   OROPKG_EXECUTION
    requires OROPKG_EXECUTION
    requires OROPKG_SUPPORT_BOOST_GRAPH
    requires OROPKG_SUPPORT_BOOST
    requires OROPKG_EXECUTION_TASK_CONTEXT

    compile VertexNode.cxx EdgeCondition.cxx
    compile FunctionGraph.cxx FunctionGraphBuilder.cxx 
    compile CommandCounter.cxx  CommandIllegal.cxx  CommandString.cxx CommandDispatch.cxx CommandExecFunction.cxx
    compile ConditionBool.cxx  ConditionBoolDataSource.cxx  ConditionBoolProperty.cxx  ConditionComposite.cxx
    compile AsynchCommandDecorator.cxx
    compile StateDescription.cxx
    compile StateMachine.cxx
    compile CommandProcessor.cxx
    compile StateMachineProcessor.cxx
    compile ProgramProcessor.cxx
    compile ProgramInterface.cxx
    compile ProgramTask.cxx StateMachineTask.cxx

    cdl_option ORONUM_EXECUTION_PROC_QUEUE_SIZE {
	display "Processor Queue Size"
	description "
The size of the command queue of the Program Processor."
	flavor data
	default_value 16
    }

}
