cdl_package OROPKG_OS {
    display "OS Abstraction Layer"
    description "
This Package groups operating system abstractions.
It defines a Thread, Mutex, IO and the capabilities
of the system for which Orocos is compiled. You
can only select one OS Package which is called the
'target'."

    include_dir rtt/os
    
    compile startstop.cxx
    compile StartStopManager.cxx
    compile Mutex.cxx
    compile ThreadInterface.cxx RunnableInterface.cxx threads.cxx
    compile PeriodicThread.cxx
    compile SingleThread.cxx
    compile main.cxx
    compile exceptions.cxx

    define_proc {
	puts $::cdl_header ""
        puts $::cdl_header "\#include <pkgconf/system.h>"
        puts $::cdl_header "\#include CYGBLD_OS_TARGET_H"
	puts $::cdl_header ""
    }

    cdl_component OROBLD_OS_EMBEDDED {
	display "Embedded Operating System"
	description "
Enable this option to run Orocos on a limited embedded
platform. This option reduces footprint and removes
C++ exceptions from the code, crippling error diagnostics. 
Leave this disabled if unsure."
	flavor bool
	default_value 0
	define ORO_EMBEDDED
	cdl_option OROBLD_OS_NOEXCEPTIONS {
	    display "Compile without exceptions (-fno-exceptions)"
	    description "
Exceptions are disabled by default during compilation. In this case,
the scripting and property marshalling packages can not
be used. Turn this option off in order to enable exceptions
and thus to allow scripting and XML marshalling."
	    default_value 1
	    define ORO_NOEXCEPTIONS
	}
    }

    cdl_option OROBLD_OS_AGNOSTIC {
	display "Hide system includes from Orocos headers."
	description "
When enabled, Orocos OS headers will not expose non standard system file
includes to the library user. In other words, every OS function call is
wrapped and they are not inlined. This makes it easier to compile
applications with Orocos headers, since no extra include paths must be
added (like /usr/realtime). Also Built-in assembly instructions
will be used instead of the system header files.
"
	flavor bool
        default_value 1
    }

    cdl_option ORONUM_OS_MAX_THREADS {
	display "The maximum number of threads in an Application."
	description "
This number is used by some buffers classes to pre-allocate per thread
data in order to allow real-time buffer operations. Most buffer
implementations have a per-buffer constructor parameter to tune this
number more precisely, meaning, to set the number of threads which 
will access a particular buffer instance concurrently.
"
	flavor data
        default_value 8
    }

    cdl_option OROCLS_OS_MINIMAL_STREAMS {
	display "Minimal streams implementation"
	description "
This provides an <iostream> like implementation of
streams, but suitable for hard realtime at the cost
of generality (so it is less configurable as the 
std C++ library). It resides in the rt_std namespace."
	flavor bool
	default_value 1
	compile rtstreams.cxx
	compile rtconversions.cxx  rtctype.cxx
    }

    cdl_option OROFUN_OS_ALTERNATE_RTTI {
	display "Alternate C++ Run Time Type Info (EXP)"
	description "
Enable to compile a C++ RTTI implementation, based on the
gcc compilers implementation. Only use if your target's
C++ libraries have no RTTI support *and* use with care.
Leave this disabled if unsure."
	flavor bool
	default_value 0
	compile rt_tinfo.cxx rt_tinfo2.cxx
	active_if OROCFG_CORELIB_EXPERIMENTAL
    }

   cdl_component OROSEM_OS_PERIODIC_THREADS_MAX_OVERRUN {
       display "Maximum number of overruns"
       description "
This option sets the maximum number of times an overrun is allowed to happen for a periodic thread.  Note that each overrun probably indicates a missed deadline.  "
       flavor data
       default_value 5
    }

    cdl_component OROPKG_OS_THREAD_SCOPE {
	display "Monitoring of Thread Execution"
	description "
When enabled, each created thread will set a bit of the 
selected port high during execution of Orocos tasks. The thread-bit
mapping is printed to the CoreLib Logger::Info stream if available.
To enable this option, enable the scope function of a device_driver component (eg the
Standard IO Ports Device Driver).
"
	flavor bool
	#calculated OROINT_DEVICE_INTERFACE_THREAD_SCOPE
	default_value 0
    }

    cdl_component OROSEM_OS_LOCK_MEMORY {
	display "Lock all virtual address space into RAM"
	description "
Enabling this option forces the OS kernel to reserve and
lock all current virtual memory in physical RAM. This guarantees
that no memory is swapped."
	flavor bool
	default_value 1
	cdl_option OROSEM_OS_LOCK_MEMORY_FUTURE {
	display "Lock future stack and heap virtual address space into RAM"
	description "
DANGER ! Enabling this option forces the OS kernel to reserve and
lock all future virtual memory in physical RAM and prevents any stack
and heap growth beyond these reserved boundaries, causing SIGSEGV if
violated. Only enable if you know what you are doing."
	flavor bool
	default_value 0
	}

    }

    # we need exactly one OS_TARGET
    cdl_interface OROINT_OS_TARGET {
	display "Target Operating System"
	flavor bool
	requires OROINT_OS_TARGET == 1
    }

    cdl_interface OROINT_OS_GLOBAL_CRT {
	display "Target calls global constructors"
	flavor bool
	requires OROINT_OS_GLOBAL_CRT <= 1
	define OS_HAVE_MANUAL_CRT
    }

    cdl_interface OROINT_OS_MAIN {
	display "Target which calls the main() function"
	flavor bool
	requires OROINT_OS_MAIN <= 1
	define OS_HAVE_MAIN
    }

    cdl_interface OROINT_OS_MAIN_THREAD {
	display "Target with MainThread class"
	flavor bool
	requires OROINT_OS_MAIN <= 1
	define OS_HAVE_MAIN_THREAD
    }

    cdl_interface OROINT_OS_LINUX_IOPERM {
	display "Support for Linux ioperm()"
	flavor bool
    }

    cdl_interface OROINT_OS_STDCXXLIB {
	display "Support for the Standard C++ Library"
	flavor bool
	implements OROINT_OS_STL_LIB
	implements OROINT_OS_STDIOSTREAM
	implements OROINT_OS_STREAMS
    }

    cdl_interface OROINT_OS_STL_LIB {
	display "Standard Template C++ Library"
	flavor bool
    }

    cdl_interface OROINT_OS_STDIOSTREAM {
	display "IO Streams (cerr,cout,...) of the Standard C++ Library"
	define HAVE_IOSTREAM
	flavor bool
    }

    cdl_interface OROINT_OS_STREAMS {
	display "Stream operations of the Standard C++ Library"
	define HAVE_STREAMS
	flavor bool
    }

    cdl_interface OROINT_OS_KERNEL {
	display "Inside-kernel interface"
	flavor bool
    }

    cdl_interface OROINT_OS_KERNEL_MODULE {
	display "Kernel module loader support"
	flavor bool
    }

    cdl_interface OROINT_OS_RECURSIVE_MUTEX {
	display "Support for recursive mutex"
	flavor bool
    }

    cdl_interface OROINT_OS_CORBA {
	display "Support for Corba."
	flavor bool
    }

    cdl_interface OROINT_OS_TAO {
	display "Support for Tao."
	flavor bool
    }
}
