
cdl_package OROPKG_EXECUTION_PROGRAM_PROCESSOR {
    display "Execution Program processing infrastructure"
    description "
A Package that provides realtime-safe program execution,
with each program statement represented by an object
which encapsulates the command to be executed."

    include_dir execution
    
    parent   OROPKG_EXECUTION
    requires OROPKG_EXECUTION
    requires OROPKG_SUPPORT_BOOST_GRAPH
    requires OROPKG_SUPPORT_BOOST
    requires OROPKG_CORELIB_STATE
    requires OROPKG_EXECUTION_TASK_CONTEXT

    compile VertexNode.cxx EdgeCondition.cxx
    compile FunctionGraph.cxx ProgramGraph.cxx 
    compile CommandCounter.cxx  CommandIllegal.cxx  CommandString.cxx  
    compile ConditionBool.cxx  ConditionBoolDataSource.cxx  ConditionBoolProperty.cxx  ConditionComposite.cxx
    compile Processor.cxx
    compile AsynchCommandDecorator.cxx
    compile StateDescription.cxx

    cdl_option ORONUM_EXECUTION_PROC_QUEUE_SIZE {
	display "Processor Queue Size"
	description "
The size of the command queue of the Program Processor."
	flavor data
	default_value 16
    }

}
