cdl_package OROPKG_DEVICE_DRIVERS_K600 {
    display "Device Drivers Real-time for Krypton K600 Measuring device"

    parent   OROPKG_DEVICE_DRIVERS

    requires OROPKG_OS_LXRT
    requires OROPKG_CORELIB_ACTIVITIES
    requires OROPKG_DEVICE_DRIVERS
    requires OROPKG_DEVICE_INTERFACE
    requires OROPKG_DEVICE_INTERFACE_IO

    include_dir rtnet
    include_files KryptonK600PositionInterfaceThread.hpp KryptonK600PositionInterfaceThread.inc
}
