

cdl_package OROPKG_OS_ECOS {
    display "OS Abstraction Layer eCos"
    description "
This package is used if you want to compile
Orocos for eCos, allowing hard
real-time userspace applications"

    include_dir os
    parent OROPKG_OS

    compile fosi.c

    implements OROINT_OS_TARGET
    implements OROINT_OS_STDCXXLIB

    requires OROPKG_SUPPORT_ECOS

}
